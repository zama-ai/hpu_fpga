// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in ksk_manager.
// ==============================================================================================

package ksk_mgr_common_cut_definition_pkg;
  localparam int KSK_CUT_NB  = 16;
endpackage
