// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
//
// // ============================================================================================== //
// // Description  : Coverage
// // ---------------------------------------------------------------------------------------------- //
// //
// // Definition of covergroups for the functional coverage of mod_reduct_barrett
// // This file is included in the module mod_reduct_barrett
// // ============================================================================================== //
// //==========================
// // Covergroups
// //==========================
// covergroup cvg_mod_reduct_barrett@(posedge clk);
//   correction : coverpoint s3_sign;
// endgroup
// //==========================
// // Covergroup creation
// //==========================
// cvg_mod_reduct_barrett cvg = new;

