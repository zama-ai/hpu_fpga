// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// /!\ Generated file. Do not modify. /!\
// Generated with ntt_gf64.sage
//
// List the PHIs for up to N=2048
// ==============================================================================================

package ntt_core_gf64_phi_phi_pkg;
  // [power of w2N]

  //========================
  // NTT forward
  //========================
  //------------------------
  // 2048
  //------------------------
  localparam [2*2048-1:0][63:0] NTT_GF64_FWD_N2048_PHI_L = {
64'hccd995a189591249,64'h88faac55bfee9b74,64'h0711cdf9749c5f45,64'hab38bf38115ea62c,
64'h112b42058dbebfae,64'h90496de5221ecc48,64'h94da9c8b77bfb9e2,64'h705cd1e9bb1779ed,
64'h4747a3d7c1b3d860,64'haef0b2d0c4ee8372,64'h0e86700baab25c06,64'h6ce8024cb0531c09,
64'h39c0852287755b1a,64'h116301356bef0471,64'hecedf13a5b40b24f,64'h80b6b6221f840fa4,
64'he6d22cc1eec41321,64'h316c0622014da8c9,64'ha318ef5c91758823,64'h47aaaec033dd535f,
64'hb688ecd818e6262f,64'hefdef1ac4cacea9d,64'h6c99fb6b94b99383,64'hbf562ae382c86418,
64'had2d79cbe38a5164,64'hc7dc8acb6bcdda91,64'h44b20bdff2803c6b,64'h3591151bb83abdfc,
64'hc7c944d72e481758,64'h3971c491d0cf36cc,64'hf99c7951df1f001f,64'h0000003fffbfffc0,
64'hedaf0561e1493bc4,64'he614a28ae8d04c3c,64'ha8b8e5b2433674d7,64'h897a64fb4f51752c,
64'hee4830fa5a03ddee,64'h0e4677cd54158713,64'hcceb51c4610f9b4a,64'h4b539e10a7c92186,
64'h76f3d90ea932c3f9,64'h8743e4862bde2b7c,64'ha9a8b348b0509d32,64'h817fb35caf13a495,
64'h94a678f8ec166100,64'hae61c7b98f42ef26,64'h815a87db60d25926,64'h585bda2e086ebc26,
64'h804f6275d269bbd0,64'hcadd83c71f60a042,64'h8614e4f8d3cae658,64'h4735f5ad465162df,
64'h0355afcd98a8e075,64'hbfeb840c3604e56a,64'h53648bc0ca776ada,64'hf9087e2b728c16ab,
64'h6f702ae179387f66,64'h4069b9747158a008,64'ha8014e1c18bf19c7,64'hc7b40bfd0e189e58,
64'h5c085176a5dae686,64'h0f4b22b2bccf84fd,64'h7309d8a2c9a00ae7,64'hdfffffff20000001,
64'hf99b32b3512b224a,64'h911f558a37fdd36f,64'h60e239bece938be9,64'h956717e6822bd4c6,
64'h4225684071b7d7f6,64'h12092dbca443d989,64'hd29b5390aef7f73d,64'h6e0b9a3cd762ef3e,
64'h08e8f47af8367b0c,64'hd5de1659589dd06f,64'h41d0ce0135564b81,64'hed9d0048b60a6382,
64'hc73810a390eeab64,64'he22c6025cd7de08f,64'h3d9dbe272b68164a,64'h9016d6c3c3f081f5,
64'hfcda45975dd88265,64'he62d80c36029b51a,64'hb4631deaf22eb105,64'h28f555d7e67baa6c,
64'h36d11d9ae31cc4c6,64'h7dfbde3529959d54,64'had933f6cd2973271,64'h17eac55c70590c83,
64'h95a5af38fc714a2d,64'hf8fb91588d79bb53,64'ha896417b5e50078e,64'h86b222a2f70757c0,
64'h18f9289ae5c902eb,64'h872e3891ba19e6da,64'h3f338f2a1be3e004,64'h00000007fff7fff8,
64'h9db5e0abbc292779,64'h9cc29450dd1a0988,64'h35171cb62866ce9b,64'h912f4c9ee9ea2ea6,
64'h5dc9061f0b407bbe,64'ha1c8cef90a82b0e3,64'hd99d6a37cc21f36a,64'h496a73c1d4f92431,
64'heede7b20f5265880,64'h90e87c90457bc570,64'hd5351668560a13a7,64'h702ff66b35e27493,
64'h1294cf1f1d82cc20,64'h55cc38f6f1e85de5,64'h502b50fb2c1a4b25,64'h4b0b7b45810dd785,
64'h1009ec4eba4d377a,64'hd95bb07823ec1409,64'h10c29c9f1a795ccb,64'h28e6beb588ca2c5c,
64'h606ab5f953151c0f,64'hd7fd7080c6c09cae,64'hca6c9177594eed5c,64'hbf210fc4ce5182d6,
64'h4dee055bef270fed,64'h080d372e8e2b1401,64'h350029c36317e339,64'h18f6817fa1c313cb,
64'h4b810a2e94bb5cd1,64'h61e96455f799f0a0,64'h2e613b143934015d,64'hfbffffff04000001,
64'hdf336655aa25644a,64'h3223eab126ffba6e,64'hec1c4736f9d2717e,64'h52ace2fc90457a99,
64'h4844ad07ce36faff,64'he24125b6b4887b32,64'h7a536a71b5defee8,64'h4dc173475aec5de8,
64'h811d1e8edf06cf62,64'h3abbc2cb0b13ba0e,64'he83a19bf46aac971,64'hddb3a00856c14c71,
64'h98e70213f21dd56d,64'h3c458c0499afbc12,64'hc7b3b7c4256d02ca,64'h7202dad8187e103f,
64'h7f9b48b28bbb104d,64'hdcc5b017ac0536a4,64'h768c63bcfe45d621,64'h851eaaba7ccf754e,
64'h46da23b31c639899,64'h8fbf7bc62532b3ab,64'hf5b267ecba52e64f,64'ha2fd58aaee0b2191,
64'h72b4b5e6bf8e2946,64'hbf1f722a71af376b,64'h5512c82f2bca00f2,64'h10d644545ee0eaf8,
64'ha31f2512bcb9205e,64'hd0e5c71177433cdc,64'h87e671e4c37c7c01,64'h00000000fffeffff,
64'hf3b6bc14978524f0,64'h1398528a1ba34131,64'ha6a2e396250cd9d4,64'h5225e9939d3d45d5,
64'h4bb920c3a1680f78,64'hb43919de8150561d,64'hdb33ad4639843e6e,64'he92d4e775a9f2487,
64'h1ddbcf641ea4cb10,64'h121d0f9208af78ae,64'h3aa6a2cceac14275,64'hae05feccc6bc4e93,
64'h025299e3e3b05984,64'h6ab9871e7e3d0bbd,64'h6a056a1f05834965,64'h69616f685021baf1,
64'hc2013d891749a6f0,64'hfb2b760e247d8282,64'ha2185393434f2b9a,64'h851cd7d63119458c,
64'h2c0d56bf0a62a382,64'h5affae0fd8d81396,64'h994d922e6b29ddac,64'h57e421f859ca305b,
64'h69bdc0ab1de4e1fe,64'he101a6e4f1c56281,64'he6a005378c62fc68,64'ha31ed02f5438627a,
64'he9702144f2976b9b,64'h0c3d2c8abef33e14,64'h65cc27622726802c,64'hff7fffff00800001,
64'hdbe66cc9f544ac8a,64'h46447d55e4dff74e,64'h5d8388e69f3a4e30,64'hea559c5eb208af54,
64'h290895a0d9c6df60,64'hdc4824b616910f67,64'h0f4a6d4e36bbdfdd,64'h09b82e68eb5d8bbd,
64'hd023a3d11be0d9ed,64'h4757785921627742,64'hfd07433708d5592f,64'hfbb674002ad8298f,
64'h731ce0421e43baae,64'hc788b17fd335f783,64'hd8f676f7c4ada05a,64'h2e405b5ae30fc208,
64'h6ff36915f177620a,64'h9b98b6027580a6d5,64'heed18c76bfc8bac5,64'h50a3d5570f99eeaa,
64'he8db4475838c7314,64'hb1f7ef7824a65676,64'h3eb64cfd774a5cca,64'hf45fab147dc16433,
64'h4e5696bc97f1c529,64'hb7e3ee44ae35e6ee,64'hcaa259052579401f,64'h021ac88a8bdc1d5f,
64'h5463e4a21797240c,64'h9a1cb8e1aee8679c,64'hf0fcce3bb86f8f81,64'h1fffffffffffe000,
64'h1e76d78292f0a49e,64'he2730a5063746827,64'h94d45c7244a19b3b,64'h6a44bd3213a7a8bb,
64'h09772418742d01ef,64'h7687233b702a0ac4,64'h5b6675a8873087ce,64'h3d25a9cecb53e491,
64'h03bb79ec83d49962,64'h4243a1f20115ef16,64'h6754d4593d58284f,64'hb5c0bfd8f8d789d3,
64'h804a533bfc760b31,64'h6d5730e36fc7a178,64'h6d40ad4380b0692d,64'hed2c2dec2a04375f,
64'h184027b122e934de,64'hdf656ec1048fb051,64'hd4430a71a869e574,64'h90a39afa462328b2,
64'hc581aad7214c5471,64'h4b5ff5c1bb1b0273,64'h9329b2454d653bb6,64'haafc843e6b39460c,
64'h4d37b81523bc9c40,64'hfc2034dbbe38ac51,64'h1cd400a6f18c5f8d,64'hd463da052a870c50,
64'hbd2e0427fe52ed74,64'h8187a590d7de67c3,64'h8cb984ebc4e4d006,64'hffefffff00100001,
64'hdb7ccd987ea89592,64'h48c88faa7c9bfeea,64'h0bb0711cd3e749c6,64'h9d4ab38b564115eb,
64'h052112b41b38dbec,64'h3b890496a2d221ed,64'h61e94da966d77bfc,64'h613705ccbd6bb178,
64'h7a047479c37c1b3e,64'hc8eaef0a642c4ee9,64'h3fa0e866c11aab26,64'h3f76ce7fe55b0532,
64'h4e639c0803c87756,64'hb8f1162f5a66bef1,64'hdb1ecede3895b40c,64'h05c80b6b5c61f841,
64'hcdfe6d21fe2eec42,64'h737316bfeeb014db,64'h7dda318e77f91759,64'hca147aaa21f33dd6,
64'h9d1b688e30718e63,64'h563efdeec494cacf,64'hc7d6c99eeee94b9a,64'hbe8bf561efb82c87,
64'he9cad2d6b2fe38a6,64'h56fc7dc855c6bcde,64'h39544b2084af2804,64'h20435911317b83ac,
64'h8a8c7c93c2f2e482,64'h9343971bb5dd0cf4,64'hfe1f99c6970df1f1,64'h03fffffffffffc00,
64'h43cedaf0125e1494,64'h3c4e6149ec6e8d05,64'hb29a8b8da8943368,64'had4897a5a274f518,
64'h212ee482ee85a03e,64'h8ed0e466ee054159,64'h4b6cceb4d0e610fa,64'he7a4b538f96a7c93,
64'hc0776f3cd07a932d,64'h4848743e0022bde3,64'h2cea9a8b07ab050a,64'hb6b817fa7f1af13b,
64'hf0094a669f8ec167,64'h0daae61c6df8f42f,64'h6da815a810160d26,64'h3da585bd654086ec,
64'h430804f5e45d269c,64'hfbecadd74091f60b,64'h9a88614db50d3caf,64'hd214735e88c46517,
64'hf8b0355a04298a8f,64'ha96bfeb79763604f,64'h5265364869aca777,64'h955f90874d6728c2,
64'h09a6f702a4779388,64'hff84069a97c7158b,64'h639a80147e318bf2,64'h1a8c7b40a550e18a,
64'h97a5c0847fca5daf,64'hb030f4b17afbccf9,64'h5197309d389c9a01,64'hfffdffff00020001,
64'hdb6f99b24fd512b3,64'hc91911f48f937fde,64'h41760e235a7ce939,64'hb3a95670cac822be,
64'h80a4225603671b7e,64'h67712092745a443e,64'h8c3d29b4acdaef80,64'h0c26e0b997ad762f,
64'h4f408e8ef86f8368,64'hf91d5de06c8589de,64'h47f41d0c98235565,64'hc7eed9cf3cab60a7,
64'h49cc7380c0790eeb,64'hf71e22c50b4cd7df,64'h9b63d9db4712b682,64'he0b9016c8b8c3f09,
64'hd9bfcda37fc5dd89,64'hae6e62d75dd6029c,64'hefbb4630eeff22ec,64'h59428f55043e67bb,
64'hb3a36d11260e31cd,64'h2ac7dfbdb892995a,64'hd8fad9331ddd2974,64'h37d17eac1df70591,
64'h5d395a5a965fc715,64'h4adf8fb8cab8d79c,64'h872a89639095e501,64'h84086b21a62f7076,
64'hd1518f91b85e5c91,64'h926872e2f6bba19f,64'hffc3f337f2e1be3f,64'h007fffffffffff80,
64'h8879db5d824bc293,64'h6789cc28dd8dd1a1,64'h16535171b512866d,64'h15a912f4b44e9ea3,
64'h4425dc901dd0b408,64'hf1da1c8bfdc0a82c,64'hc96d99d5da1cc220,64'hbcf496a67f2d4f93,
64'h780eede73a0f5266,64'ha9090e87200457bd,64'hc59d5350a0f560a2,64'hb6d702feafe35e28,
64'h3e01294cb3f1d82d,64'h21b55cc36dbf1e86,64'h4db502b4c202c1a5,64'h87b4b0b72ca810de,
64'h8861009e3c8ba4d4,64'hbf7d95ba48123ec2,64'h33510c2996a1a796,64'h3a428e6bb1188ca3,
64'h3f1606ab20853152,64'h352d7fd6d2ec6c0a,64'h2a4ca6c8ed3594ef,64'hd2abf21029ace519,
64'h0134dee0548ef271,64'hbff080d2b2f8e2b2,64'hcc735001cfc6317f,64'hc3518f6754aa1c32,
64'h32f4b8106ff94bb6,64'hf6061e954f5f79a0,64'hea32e612c7139341,64'hffffbfff00004001,
64'hbb6df335a9faa257,64'h5923223e51f26ffc,64'he82ec1c38b4f9d28,64'h56752acdd9590458,
64'h5014844a806ce370,64'h4cee24120e8b4888,64'h1187a536959b5df0,64'h2184dc1712f5aec6,
64'h09e811d1df0df06d,64'h5f23abbbcd90b13c,64'h68fe83a133046aad,64'h38fddb39c7956c15,
64'ha9398e6f780f21de,64'h3ee3c45881699afc,64'hd36c7b3aa8e256d1,64'hfc17202cb17187e2,
64'hfb37f9b38ff8bbb2,64'h95cdcc5a6bbac054,64'h9df768c59ddfe45e,64'hab2851ea0087ccf8,
64'h76746da1c4c1c63a,64'hc558fbf6f712532c,64'h9b1f5b25e3bba52f,64'he6fa2fd4a3bee0b3,
64'h6ba72b4af2cbf8e3,64'h895bf1f699571af4,64'hf0e5512b9212bca1,64'h50810d63f4c5ee0f,
64'hfa2a31f1570bcb93,64'h324d0e5c3ed77434,64'h3ff87e66de5c37c8,64'h000ffffffffffff0,
64'hb10f3b6b10497853,64'hecf139843bb1ba35,64'h62ca6a2dd6a250ce,64'ha2b5225df689d3d5,
64'h0884bb9203ba1681,64'h9e3b4390ffb81506,64'h192db33abb439844,64'hb79e92d42fe5a9f3,
64'h4f01ddbca741ea4d,64'h752121d084008af8,64'hd8b3aa69541eac15,64'h16dae05fd5fc6bc5,
64'h67c02529367e3b06,64'h4436ab982db7e3d1,64'h69b6a05638405835,64'h50f69616a595021c,
64'h910c20134791749b,64'hd7efb2b6890247d9,64'h466a2184f2d434f3,64'ha74851ccd6231195,
64'hc7e2c0d4a410a62b,64'hc6a5affa1a5d8d82,64'h254994d8fda6b29e,64'hfa557e4125359ca4,
64'he0269bdb2a91de4f,64'hd7fe1019965f1c57,64'h398e6a0019f8c630,64'hd86a31ec2a954387,
64'h465e9701cdff2977,64'h1ec0c3d2a9ebef34,64'hfd465cc178e27269,64'hfffff7ff00000801,
64'h376dbe66953f544b,64'h8b2464474a3e4e00,64'h1d05d8387169f3a5,64'h0acea559bb2b208b,
64'h0a029089500d9c6e,64'h099dc48241d16911,64'h0230f4a6d2b36bbe,64'h44309b82a25eb5d9,
64'h613d0239dbe1be0e,64'h8be47576f9b21628,64'h6d1fd073c6608d56,64'h671fbb66d8f2ad83,
64'h552731cdaf01e43c,64'h87dc788a902d3360,64'hfa6d8f66751c4adb,64'hdf82e404d62e30fd,
64'hdf66ff35b1ff1777,64'h92b9b98acd77580b,64'h53beed1873bbfc8c,64'h15650a3d4010f99f,
64'hcece8db3789838c8,64'h98ab1f7e5ee24a66,64'h3363eb649c7774a6,64'hbcdf45f9f477dc17,
64'had74e568be597f1d,64'h912b7e3e532ae35f,64'hfe1caa2492425795,64'h2a1021ac5e98bdc2,
64'hbf45463d8ae17973,64'h8649a1cb07daee87,64'h07ff0fccdbcb86f9,64'h0001fffffffffffe,
64'hb621e76cc2092f0b,64'h7d9e273027763747,64'h4c594d457ad44a1a,64'h7456a44b5ed13a7b,
64'he1109771607742d1,64'h53c76871dff702a1,64'h8325b666d7687309,64'hb6f3d259e5fcb53f,
64'h69e03bb734e83d4a,64'h0ea4243a1080115f,64'h7b16754cca83d583,64'h62db5c0b9abf8d79,
64'h4cf804a4e6cfc761,64'he886d57225b6fc7b,64'h6d36d40a67080b07,64'h8a1ed2c254b2a044,
64'hb2218401c8f22e94,64'hfafdf655f12048fc,64'ha8cd442ffe5a869f,64'h74e90a393ac46233,
64'hb8fc5819f48214c6,64'hd8d4b5fe834bb1b1,64'h44a9329adfb4d654,64'h9f4aafc7a4a6b395,
64'h3c04d37b45523bca,64'h3affc20312cbe38b,64'h0731cd40033f18c6,64'h3b0d463d6552a871,
64'h28cbd2e019bfe52f,64'h83d81879d53d7de7,64'hffa8cb974f1c4e4e,64'hfffffeff00000101,
64'ha6edb7cc32a7ea8a,64'h11648c88e947c9c0,64'h63a0bb06ae2d3e75,64'ha159d4aa97656412,
64'h41405210ea01b38e,64'he133b88f683a2d23,64'h40461e949a566d78,64'he886136f744bd6bc,
64'h4c27a046fb7c37c2,64'h117c8eaedf3642c5,64'h4da3fa0e38cc11ab,64'hace3f76c3b1e55b1,
64'h8aa4e63935e03c88,64'h10fb8f115205a66c,64'hbf4db1ec2ea3895c,64'h7bf05c803ac5c620,
64'h3becdfe6963fe2ef,64'hb2573730b9aeeb02,64'h8a77dda28e777f92,64'h22aca14788021f34,
64'h19d9d1b66f130719,64'h531563ef8bdc494d,64'h466c7d6c538eee95,64'h379be8bf1e8efb83,
64'h75ae9cacb7cb2fe4,64'h32256fc7aa655c6c,64'h7fc3954432484af3,64'hc5420434cbd317b9,
64'hb7e8a8c7115c2f2f,64'h30c9343940fb5dd1,64'he0ffe1f8bb7970e0,64'h40003fffc0000000,
64'hb6c43cecf84125e2,64'h2fb3c4e5e4eec6e9,64'hc98b29a7ef5a8944,64'hae8ad488cbda2750,
64'hfc2212ed4c0ee85b,64'hea78ed0d5bfee055,64'hf064b6cbfaed0e62,64'h36de7a4b1cbf96a8,
64'hcd3c0776269d07aa,64'h21d484872210022c,64'haf62cea8f9507ab1,64'hec5b6b809357f1b0,
64'he99f0093bcd9f8ed,64'hbd10daada4b6df90,64'h2da6da812ce10161,64'h9143da57ca965409,
64'h9644307fb91e45d3,64'h9f5fbeca3e240920,64'h3519a885dfcb50d4,64'hae9d214687588c47,
64'h571f8b02fe904299,64'hfb1a96bef0697637,64'h88952652dbf69acb,64'h73e955f89494d673,
64'hc7809a6ea8aa477a,64'ha75ff83fc2597c72,64'h40e639a7c067e319,64'he761a8c6ccaa550f,
64'h25197a5be337fca6,64'h307b030f1aa7afbd,64'h5ff51972a9e389ca,64'hffffffdf00000021,
64'hd4ddb6f8c654fd52,64'h022c91911d28f938,64'h6c74176075c5a7cf,64'hd42b3a9492ecac83,
64'h48280a41dd403672,64'hbc2677114d0745a5,64'h0808c3d2934acdaf,64'h9d10c26d6e897ad8,
64'hc984f4081f6f86f9,64'h622f91d57be6c859,64'ha9b47f4127198236,64'hf59c7eeca763cab7,
64'h11549cc726bc0791,64'h821f71e1aa40b4ce,64'h97e9b63d05d4712c,64'h0f7e0b900758b8c4,
64'h277d9bfcb2c7fc5e,64'hd64ae6e55735dd61,64'hd14efbb391ceeff3,64'h84559428710043e7,
64'he33b3a35ede260e4,64'h6a62ac7d917b892a,64'h68cd8fad2a71ddd3,64'ha6f37d1743d1df71,
64'h8eb5d39516f965fd,64'h8644adf8754cab8e,64'haff872a7e649095f,64'hf8a84085b97a62f8,
64'h36fd1518c22b85e6,64'he6192686481f6bbb,64'h1c1ffc3f176f2e1c,64'h080007fff8000000,
64'hd6d8879cdf0824bd,64'he5f6789bdc9dd8de,64'h993165347deb5129,64'h15d15a91197b44ea,
64'hbf84425d0981dd0c,64'h7d4f1da14b7fdc0b,64'hde0c96d8bf5da1cd,64'h06dbcf496397f2d5,
64'hd9a780ee04d3a0f6,64'h843a909064420046,64'hf5ec59d43f2a0f57,64'h1d8b6d70126afe36,
64'h7d33e012179b3f1e,64'h17a21b55b496dbf2,64'he5b4db4f459c202d,64'hf2287b4a1952ca82,
64'hb2c8860f5723c8bb,64'h13ebf7d947c48124,64'h86a335103bf96a1b,64'h35d3a428b0eb1189,
64'heae3f15f7fd20854,64'h3f6352d7be0d2ec7,64'hb112a4c9bb7ed35a,64'hae7d2abe72929acf,
64'hd8f0134d151548f0,64'hd4ebff07384b2f8f,64'he81cc734180cfc64,64'h3cec3518b9954aa2,
64'h44a32f4b3c66ff95,64'h660f60618354f5f8,64'hcbfea32d953c713a,64'hfffffffb00000005,
64'hda9bb6de58ca9fab,64'h0045923223a51f27,64'h2d8e82ebeeb8b4fa,64'hba856751f25d9591,
64'hc90501477ba806cf,64'h7784cee1c9a0e8b5,64'h2101187a326959b6,64'h13a2184dadd12f5b,
64'hf9309e8023edf0e0,64'hec45f239cf7cd90c,64'h55368fe7e4e33047,64'h3eb38fdd74ec7957,
64'he22a939804d780f3,64'h5043ee3bf548169a,64'h92fd36c720ba8e26,64'h81efc17180eb1719,
64'h44efb37f5658ff8c,64'hfac95cdbcae6bbad,64'hba29df75d239ddff,64'h308ab284ee20087d,
64'h9c6767463dbc4c1d,64'hcd4c558ef22f7126,64'had19b1f5054e3bbb,64'hf4de6fa2087a3bef,
64'h71d6ba7242df2cc0,64'h50c895becea99572,64'h35ff0e54dcc9212c,64'h1f150810b72f4c5f,
64'h46dfa2a2d84570bd,64'hbcc324d02903ed78,64'h8383ff8762ede5c4,64'h010000ffff000000,
64'h7adb10f33be10498,64'h5cbecf133b93bb1c,64'hf3262ca5afbd6a26,64'hc2ba2b51632f689e,
64'h97f0884b21303ba2,64'hafa9e3b3896ffb82,64'h7bc192dab7ebb43a,64'h60db79e8cc72fe5b,
64'h5b34f01d809a741f,64'h50875211cc884009,64'h3ebd8b3a67e541eb,64'h43b16dadc24d5fc7,
64'h4fa67c0202f367e4,64'hc2f44369f692db7f,64'h7cb69b6988b38406,64'hde450f68832a5951,
64'hb65910c14ae47918,64'h827d7efaa8f89025,64'hb0d466a1677f2d44,64'he6ba7484361d6232,
64'h9d5c7e2b6ffa410b,64'h27ec6a5ad7c1a5d9,64'hd6225498776fda6c,64'h35cfa557ae52535a,
64'h1b1e0269a2a2a91e,64'h3a9d7fe0c70965f2,64'h9d0398e603019f8d,64'hc79d86a25732a955,
64'h689465e9078cdff3,64'h0cc1ec0c306a9ebf,64'hd97fd464f2a78e28,64'h7fffffff00000001,
64'hbb5376db2b1953f6,64'h2008b2462474a3e5,64'hc5b1d05cbdd716a0,64'hf750ace95e4bb2b3,
64'h3920a028cf7500da,64'h6ef099dbd9341d17,64'h4420230f064d2b37,64'ha274430915ba25ec,
64'h1f2613d0047dbe1c,64'h9d88be46b9ef9b22,64'h2aa6d1fcdc9c6609,64'h27d671fb8e9d8f2b,
64'hbc455272609af01f,64'hca087dc6bea902d4,64'h525fa6d8a41751c5,64'hf03df82d501d62e4,
64'h889df66f6acb1ff2,64'h7f592b9b195cd776,64'h37453bee9a473bc0,64'h661156503dc40110,
64'h738cece867b78984,64'h59a98ab19e45ee25,64'hb5a3363e00a9c778,64'h3e9bcdf4210f477e,
64'h0e3ad74e485be598,64'hca1912b719d532af,64'h86bfe1ca1b992426,64'h23e2a101f6e5e98c,
64'h68dbf453fb08ae18,64'h1798649a05207daf,64'h90707ff06c5dbcb9,64'h0020001fffe00000,
64'h0f5b621e677c2093,64'h8b97d9e1e7727764,64'h5e64c59475f7ad45,64'h58574569ec65ed14,
64'hd2fe1108a4260775,64'hd5f53c75b12dff71,64'hcf78325a96fd7688,64'hac1b6f3c798e5fcc,
64'h2b669e0390134e84,64'hea10ea4159910802,64'ha7d7b166acfca83e,64'h28762db59849abf9,
64'h89f4cf7fc05e6cfd,64'h385e886d1ed25b70,64'h4f96d36cf1167081,64'hfbc8a1ec30654b2b,
64'h16cb2218295c8f23,64'h704fafdef51f1205,64'h961a8cd3acefe5a9,64'hdcd74e8fc6c3ac47,
64'hb3ab8fc4cdff4822,64'he4fd8d4a7af834bc,64'h9ac44a928eedfb4e,64'hc6b9f4aa35ca4a6c,
64'h4363c04cf4545524,64'hc753affb58e12cbf,64'h73a0731c606033f2,64'h78f3b0d3eae6552b,
64'had128cbc80f19bff,64'h21983d81660d53d8,64'h1b2ffa8c9e54f1c5,64'hefffffff00000001,
64'h576a6edb25632a7f,64'h64011648648e947d,64'h18b63a0b97bae2d4,64'hbeea159c8bc97657,
64'hc724140459eea01c,64'h2dde133b5b2683a3,64'h28840461c0c9a567,64'h944e8860a2b744be,
64'h83e4c279808fb7c4,64'hd3b117c8173df365,64'he554da3ebb938cc2,64'ha4face3ed1d3b1e6,
64'h3788aa4e2c135e04,64'h99410fb857d5205b,64'h6a4bf4dab482ea39,64'h9e07bf052a03ac5d,
64'hd113becd2d5963ff,64'h4feb2573232b9aef,64'h06e8a77dd348e778,64'h0cc22aca07b88022,
64'h8e719d9c8cf6f131,64'h6b353155d3c8bdc5,64'h16b466c7c01538ef,64'h47d379be4421e8f0,
64'h01c75ae9c90b7cb3,64'h39432256c33aa656,64'h50d7fc3903732485,64'h847c541fbedcbd32,
64'h0d1b7e8a7f6115c3,64'h22f30c9320a40fb6,64'hf20e0ffd2d8bb798,64'h00040003fffc0000,
64'ha1eb6c432cef8413,64'h9172fb3bbcee4eed,64'h6bcc98b22ebef5a9,64'h8b0ae8acbd8cbda3,
64'h7a5fc220b484c0ef,64'hfabea78dd625bfef,64'h19ef064b52dfaed1,64'h95836de70f31cbfa,
64'h856cd3bff20269d1,64'hdd421d476b322101,64'h54faf62c959f9508,64'he50ec5b5d3093580,
64'h713e99ef980bcda0,64'h070bd10da3da4b6e,64'he9f2da6cbe22ce11,64'hbf79143ce60ca966,
64'ha2d96442652b91e5,64'h6e09f5fb7ea3e241,64'hf2c35199959dfcb6,64'h3b9ae9d1d8d87589,
64'hd67571f7d9bfe905,64'h9c9fb1a8cf5f0698,64'h5358895211ddbf6a,64'h98d73e94c6b9494e,
64'h886c78091e8a8aa5,64'h38ea75ff4b1c2598,64'hce740e62cc0c067f,64'haf1e7619dd5ccaa6,
64'h35a25197701e3380,64'h043307b02cc1aa7b,64'h6365ff5133ca9e39,64'hfdffffff00000001,
64'h2aed4ddb44ac6550,64'h6c8022c8ac91d290,64'h8316c740f2f75c5b,64'h37dd42b371792ecb,
64'h98e482800b3dd404,64'ha5bbc266cb64d075,64'h2510808c181934ad,64'h5289d10bd456e898,
64'h907c984eb011f6f9,64'h7a7622f8a2e7be6d,64'hdcaa9b4717727199,64'h549f59c79a3a763d,
64'h86f1154945826bc1,64'hb32821f66afaa40c,64'hed497e9a76905d48,64'h73c0f7e04540758c,
64'h3a2277d985ab2c80,64'h29fd64ae4465735e,64'h00dd14efba691cef,64'hc198455880f71005,
64'hf1ce33b2b19ede27,64'h6d66a62a5a7917b9,64'h22d68cd8d802a71e,64'h08fa6f37c8843d1e,
64'ha038eb5c99216f97,64'h4728644a986754cb,64'h6a1aff86c06e6491,64'hd08f8a8337db97a7,
64'ha1a36fd0afec22b9,64'h445e6192241481f7,64'h1e41c1ffa5b176f3,64'h000080007fff8000,
64'hb43d6d87c59df083,64'h722e5f67179dc9de,64'hed79931565d7deb6,64'hb1615d14f7b197b5,
64'h2f4bf843f690981e,64'h3f57d4f19ac4b7fe,64'he33de0c88a5bf5db,64'hd2b06dbc21e63980,
64'hf0ad9a771e404d3b,64'hfba843a80d664421,64'h0a9f5ec592b3f2a1,64'h1ca1d8b6ba6126b0,
64'h0e27d33df30179b4,64'h40e17a21747b496e,64'hfd3e5b4cb7c459c3,64'h57ef22875cc1952d,
64'h745b2c87eca5723d,64'hedc13ebe8fd47c49,64'h5e586a32f2b3bf97,64'he7735d395b1b0eb2,
64'h7aceae3e9b37fd21,64'h1393f63519ebe0d3,64'hca6b1129823bb7ee,64'h531ae7d258d7292a,
64'h710d8f00c3d15155,64'h071d4ebfe96384b3,64'h39ce81cc398180d0,64'h55e3cec2fbab9955,
64'h06b44a32ee03c670,64'ha08660f565983550,64'hec6cbfe9467953c8,64'hffbfffff00000001,
64'h055da9bb68958caa,64'h0d90045915923a52,64'hb062d8e77e5eeb8c,64'ha6fba855ce2f25da,
64'h931c904f8167ba81,64'h74b7784c796c9a0f,64'h64a2101123032696,64'h0a513a217a8add13,
64'hf20f9308f6023ee0,64'h6f4ec45eb45cf7ce,64'hfb95536802ee4e34,64'h6a93eb3893474ec8,
64'hf0de22a848b04d79,64'h9665043e4d5f5482,64'h1da92fd34ed20ba9,64'h8e781efb88a80eb2,
64'h07444efb30b56590,64'h453fac95888cae6c,64'h201ba29dd74d239e,64'h783308aab01ee201,
64'h3e39c6763633dbc5,64'hedacd4c46b4f22f8,64'h445ad19adb0054e4,64'h411f4de6b91087a4,
64'h34071d6b73242df3,64'ha8e50c88b30cea9a,64'hed435feff80dcc93,64'h3a11f15046fb72f5,
64'hf4346df935fd8458,64'h288bcc322482903f,64'ha3c8383f54b62edf,64'h000010000ffff000,
64'hb687adb058b3be11,64'h4e45cbeca2f3b93c,64'h5daf32626cbafbd7,64'h762c2ba23ef632f7,
64'h45e97f083ed21304,64'h47eafa9df3589700,64'hbc67bc18714b7ebc,64'h1a560db7843cc730,
64'hbe15b34e43c809a8,64'hff75087421acc885,64'he153ebd7d2567e55,64'h03943b16d74c24d6,
64'h81c4fa673e602f37,64'h481c2f43ee8f692e,64'hbfa7cb68f6f88b39,64'h6afde4508b9832a6,
64'h6e8b65909d94ae48,64'hfdb827d6f1fa8f8a,64'h2bcb0d463e5677f3,64'hdcee6ba66b6361d7,
64'hef59d5c6f366ffa5,64'ha2727ec6033d7c1b,64'h594d6224f04776fe,64'hca635cf98b1ae526,
64'h6e21b1dfb87a2a2b,64'ha0e3a9d75d2c7097,64'h0739d0398730301a,64'h6abc79d7ff75732b,
64'h00d689465dc078ce,64'h1410cc1eacb306aa,64'h1d8d97fd28cf2a79,64'hfff7ffff00000001,
64'hc0abb536ad12b196,64'hc1b2008a62b2474b,64'h960c5b1c6fcbdd72,64'hd4df7509f9c5e4bc,
64'hf2639209102cf751,64'h2e96ef096f2d9342,64'h4c944201e46064d3,64'ha14a27438f515ba3,
64'h1e41f2611ec047dc,64'h4de9d88b968b9efa,64'h9f72aa6c805dc9c7,64'h0d527d671268e9d9,
64'hfe1bc454291609b0,64'hd2cca08709abea91,64'he3b525f989da4176,64'hd1cf03deb11501d7,
64'h00e889df6616acb2,64'h88a7f592311195ce,64'h440374537ae9a474,64'hef0661147603dc41,
64'h67c738ce66c67b79,64'h1db59a988d69e45f,64'h888b5a32db600a9d,64'h8823e9bc572210f5,
64'ha680e3acce6485bf,64'hd51ca19056619d54,64'hbda86bfd5f01b993,64'h67423e29a8df6e5f,
64'h1e868dbf26bfb08b,64'h2511798624905208,64'h34790707ca96c5dc,64'h0000020001fffe00,
64'hf6d0f5b52b1677c3,64'h89c8b97d145e7728,64'h2bb5e64c2d975f7b,64'h2ec5857427dec65f,
64'h88bd2fe087da4261,64'h08fd5f53be6b12e0,64'h978cf7828e296fd8,64'h034ac1b6f08798e6,
64'h17c2b669c8790135,64'h7feea10e24359911,64'h7c2a7d7a9a4acfcb,64'h407287629ae9849b,
64'h30389f4cc7cc05e7,64'h490385e83dd1ed26,64'hf7f4f96c3edf1168,64'h4d5fbc89d1730655,
64'h0dd16cb213b295c9,64'hdfb704fa1e3f51f2,64'ha57961a827caceff,64'h3b9dcd74ad6c6c3b,
64'h7deb3ab87e6cdff5,64'hb44e4fd82067af84,64'h4b29ac445e08eee0,64'h594c6b9ef1635ca5,
64'hadc4363b570f4546,64'h341c753acba58e13,64'hc0e73a0670e60604,64'had578f3a5feeae66,
64'h401ad1288bb80f1a,64'hc2821983159660d6,64'he3b1b2fec519e550,64'hfffeffff00000001,
64'h581576a695a25633,64'hb8364010ac5648ea,64'hd2c18b62cdf97baf,64'h9a9beea0bf38bc98,
64'hfe4c724042059eeb,64'hc5d2dde06de5b269,64'ha992883f9c8c0c9b,64'hb42944e7d1ea2b75,
64'h83c83e4ba3d808fc,64'hc9bd3b10b2d173e0,64'h33ee554d700bb939,64'he1aa4fac024d1d3c,
64'h1fc3788a8522c136,64'hfa59941001357d53,64'h5c76a4bef13b482f,64'h3a39e07bb622a03b,
64'hc01d113b2cc2d597,64'h5114feb2062232ba,64'h88806e89ef5d348f,64'hfde0cc21aec07b89,
64'hecf8e718ecd8cf70,64'h23b6b352f1ad3c8c,64'h71116b45fb6c0154,64'h71047d372ae4421f,
64'h34d01c7579cc90b8,64'h9aa394318acc33ab,64'hb7b50d7f0be03733,64'h2ce847c5151bedcc,
64'ha3d0d1b744d7f612,64'h04a22f30c4920a41,64'h868f20e07952d8bc,64'h00000040003fffc0,
64'hbeda1eb60562cef9,64'h1139172fa28bcee5,64'ha576bcc8e5b2ebf0,64'h25d8b0ae64fbd8cc,
64'hf117a5fb30fb484d,64'h011fabea77cd625c,64'h12f19ef051c52dfb,64'h406958369e10f31d,
64'h62f856ccd90f2027,64'heffdd420e486b323,64'haf854faeb34959fa,64'ha80e50ebb35d3094,
64'h260713e978f980bd,64'h492070bcc7ba3da5,64'h1efe9f2d87dbe22d,64'h69abf790da2e60cb,
64'he1ba2d95627652ba,64'hdbf6e09e83c7ea3f,64'h34af2c34e4f959e0,64'ha773b9adf5ad8d88,
64'h6fbd6756afcd9bff,64'h9689c9fa840cf5f1,64'h096535888bc11ddc,64'h6b298d737e2c6b95,
64'h55b886c72ae1e8a9,64'ha6838ea6b974b1c3,64'h981ce7404e1cc0c1,64'h55aaf1e70bfdd5cd,
64'hc8035a24517701e4,64'h5850433022b2cc1b,64'h1c76365fd8a33caa,64'hffffdfff00000001,
64'hab02aed432b44ac7,64'hd706c801558ac91e,64'h3a58316c39bf2f76,64'h13537dd417e71793,
64'hbfc98e476840b3de,64'hf8ba5bbb2dbcb64e,64'hb532510753918194,64'h7685289c9a3d456f,
64'h907907c8f47b0120,64'h1937a762165a2e7c,64'he67dcaa8ce017728,64'h9c3549f50049a3a8,
64'h43f86f1110a45827,64'hbf4b32816026afab,64'h2b8ed497be276906,64'ha7473c0ed6c45408,
64'h3803a22745985ab3,64'hca229fd580c44658,64'h31100dd11deba692,64'hffbc198355d80f72,
64'h1d9f1ce31d9b19ee,64'h8476d669de35a792,64'h8e222d683f6d802b,64'h2e208fa6c55c8844,
64'h069a038eaf399217,64'hb354728591598676,64'hb6f6a1af417c06e7,64'h859d08f822a37dba,
64'hd47a1a36289afec3,64'he09445e538924149,64'h90d1e41b8f2a5b18,64'h000000080007fff8,
64'hf7db43d5e0ac59e0,64'h622722e5945179dd,64'h14aed7991cb65d7e,64'h84bb16154c9f7b1a,
64'h7e22f4bf061f690a,64'h8023f57ccef9ac4c,64'ha25e33dd6a38a5c0,64'h680d2b0673c21e64,
64'h2c5f0ad97b21e405,64'hbdffba837c90d665,64'hd5f0a9f516692b40,64'h9501ca1cf66ba613,
64'h64c0e27ccf1f3018,64'h69240e1738f747b5,64'h63dfd3e550fb7c46,64'had357ef17b45cc1a,
64'hdc3745b1ec4eca58,64'h3b7edc13b078fd48,64'h0695e5869c9f2b3c,64'h14ee7735beb5b1b1,
64'h2df7aceab5f9b380,64'hf2d1393e70819ebf,64'h812ca6b0917823bc,64'h6d6531ae0fc58d73,
64'heab710d8055c3d16,64'hb4d071d4372e9639,64'hf3039ce729c39819,64'h6ab55e3c817fbaba,
64'h99006b440a2ee03d,64'hab0a086564565984,64'hc38ec6cb3b146796,64'hfffffbff00000001,
64'h356055da66568959,64'h5ae0d8ffeab15924,64'h474b062d4737e5ef,64'ha26a6fb9e2fce2f3,
64'h57f931c8ad08167c,64'h5f174b7725b796ca,64'h96a64a206a723033,64'h2ed0a5137347a8ae,
64'h120f20f91e8f6024,64'h8326f4ebc2cb45d0,64'h1ccfb95519c02ee5,64'h1386a93ea0093475,
64'h287f0de202148b05,64'hb7e9664f8c04d5f6,64'h4571da92b7c4ed21,64'h14e8e781dad88a81,
64'ha700744448b30b57,64'h194453fab01888cb,64'hc62201b963bd74d3,64'hdff7832faabb01ef,
64'h43b3e39c23b3633e,64'hd08edacc7bc6b4f3,64'hb1c445ac67edb006,64'h85c411f458ab9109,
64'h20d34071b5e73243,64'h566a8e50722b30cf,64'h36ded435c82f80dd,64'hd0b3a11e44546fb8,
64'hba8f434625135fd9,64'hfc1288bbc712482a,64'h121a3c8371e54b63,64'h000000010000ffff,
64'h1efb687abc158b3c,64'h6c44e45c528a2f3c,64'h4295daf2e396cbb0,64'hd09762c1e993ef64,
64'hcfc45e9720c3ed22,64'h90047eaf19df358a,64'h144bc67bad4714b8,64'h8d01a5604e7843cd,
64'h658be15acf643c81,64'h77bff7500f921acd,64'h1abe153ea2cd2568,64'hb2a03942fecd74c3,
64'h0c981c4f99e3e603,64'h6d2481c2871ee8f7,64'h4c7bfa7c6a1f6f89,64'hd5a6afdd6f68b984,
64'h1b86e8b63d89d94b,64'h076fdb82760f1fa9,64'h80d2bcb05393e568,64'he29dcee5d7d6b637,
64'h05bef59d56bf3670,64'h3e5a2727ae1033d8,64'h902594d5922f0478,64'hadaca63521f8b1af,
64'h5d56e21ac0ab87a3,64'hf69a0e39a6e5d2c8,64'hfe60739c05387304,64'hcd56abc6d02ff758,
64'h73200d682145dc08,64'h9561410c2c8acb31,64'h5871d8d927628cf3,64'hffffff7f00000001,
64'he6ac0aba6ccad12c,64'h8b5c1b1f7d562b25,64'h28e960c588e6fcbe,64'hb44d4df69c5f9c5f,
64'h8aff263895a102d0,64'hcbe2e96e24b6f2da,64'hb2d4c9436d4e4607,64'h45da14a22e68f516,
64'h8241e41ea3d1ec05,64'h1064de9d785968ba,64'h6399f72a433805dd,64'h6270d5277401268f,
64'h650fe1bbe0429161,64'h56fd2cc9b1809abf,64'he8ae3b5176f89da5,64'he29d1cef5b5b1151,
64'h34e00e886916616b,64'ha3288a7eb603111a,64'hb8c440368c77ae9b,64'h3bfef065d557603e,
64'h48767c7344766c68,64'hba11db58ef78d69f,64'h563888b54cfdb601,64'hf0b8823dab157222,
64'ha41a680d96bce649,64'h2acd51c9ee45661a,64'h66dbda865905f01c,64'h1a167423c88a8df7,
64'hf751e867e4a26bfc,64'hdf825116b8e24906,64'ha243478fce3ca96d,64'h2000000000002000,
64'h83df6d0ed782b168,64'h8d889c8b0a5145e8,64'h0852bb5e5c72d976,64'h9a12ec57bd327ded,
64'hd9f88bd224187da5,64'hd2008fd5233be6b2,64'h028978cf75a8e297,64'h71a034aba9cf087a,
64'hecb17c2a79ec8791,64'h6ef7fee9a1f2435a,64'h0357c2a7d459a4ad,64'hb6540727bfd9ae99,
64'ha1930389533c7cc1,64'h2da4903830e3dd1f,64'he98f7f4ead43edf2,64'h9ab4d5fb2ded1731,
64'ha370dd1627b13b2a,64'he0edfb6f6ec1e3f6,64'h101a57960a727cad,64'h3c53b9dc9afad6c7,
64'h00b7deb3aad7e6ce,64'h07cb44e4f5c2067b,64'h1204b29ab245e08f,64'h35b594c6843f1636,
64'habaadc42b81570f5,64'h1ed341c734dcba59,64'h9fcc0e7300a70e61,64'h19aad578da05feeb,
64'h0e6401ad0428bb81,64'hf2ac2820a5915967,64'hab0e3b1a84ec519f,64'hffffffef00000001,
64'h9cd58156cd995a26,64'h716b83638faac565,64'h451d2c18711cdf98,64'h3689a9beb38bf38c,
64'h115fe4c712b4205a,64'hd97c5d2d0496de5c,64'h365a99284da9c8c1,64'h48bb429405cd1ea3,
64'h70483c83747a3d81,64'hc20c9bd2ef0b2d18,64'h6c733ee4e86700bc,64'h2c4e1aa4ce8024d2,
64'heca1fc369c08522d,64'h2adfa59916301358,64'h7d15c769cedf13b5,64'hfc53a39d0b6b622b,
64'ha69c01d06d22cc2e,64'hd465114f16c06224,64'hb7188806318ef5d4,64'h477fde0c7aaaec08,
64'h090ecf8e688ecd8d,64'h37423b6afdef1ad4,64'heac71115c99fb6c1,64'hde171046f562ae45,
64'hf4834d00d2d79cca,64'hc559aa387dc8acc4,64'h8cdb7b504b20be04,64'h2342ce84591151bf,
64'h9eea3d0c7c944d80,64'h5bf04a22971c4921,64'h744868f199c7952e,64'h0400000000000400,
64'h107beda1daf0562d,64'h11b11391614a28bd,64'h410a576b8b8e5b2f,64'h73425d8a97a64fbe,
64'h7b3f1179e4830fb5,64'hda4011f9e4677cd7,64'h20512f19ceb51c53,64'hce340694b539e110,
64'hfd962f846f3d90f3,64'hcddeffdc743e486c,64'h606af8549a8b3496,64'hf6ca80e417fb35d4,
64'hf43260704a678f99,64'h25b49206e61c7ba4,64'hdd31efe915a87dbf,64'hf3569abe85bda2e7,
64'hd46e1ba204f62766,64'h5c1dbf6dadd83c7f,64'h62034af2614e4f96,64'h278a773b735f5ad9,
64'h4016fbd6355afcda,64'ha0f9689bfeb840d0,64'h224096533648bc12,64'h46b6b2989087e2c7,
64'h75755b87f702ae1f,64'he3da6838069b974c,64'hf3f981cd8014e1cd,64'ha3355aae7b40bfde,
64'he1cc8034c0851771,64'h3e558503f4b22b2d,64'h3561c763309d8a34,64'hfffffffd00000001,
64'h539ab02a99b32b45,64'h6e2d706c11f558ad,64'h08a3a5830e239bf3,64'h86d1353756717e72,
64'hc22bfc982256840c,64'h9b2f8ba52092dbcc,64'he6cb532429b53919,64'ha9176851e0b9a3d5,
64'hee09078f8e8f47b1,64'h1841937a5de165a3,64'h8d8e67dc1d0ce018,64'hc589c353d9d0049b,
64'h7d943f8673810a46,64'h055bf4b322c6026b,64'h6fa2b8ecd9dbe277,64'hbf8a7473016d6c46,
64'h54d38039cda45986,64'h9a8ca22962d80c45,64'h96e311004631debb,64'h08effbc18f555d81,
64'h6121d9f16d11d9b2,64'h86e8476cdfbde35b,64'hfd58e221d933f6d9,64'h7bc2e2087eac55c9,
64'hde90699f5a5af39a,64'h98ab35468fb91599,64'h919b6f69896417c1,64'h246859d06b222a38,
64'h13dd47a18f9289b0,64'heb7e094372e38925,64'h4e890d1df338f2a6,64'h0080000000000080,
64'h620f7db3db5e0ac6,64'h62362271cc294518,64'h28214aed5171cb66,64'h4e684bb112f4c9f8,
64'h6f67e22edc9061f7,64'h3b48023f1c8cef9b,64'ha40a25e299d6a38b,64'h19c680d296a73c22,
64'hbfb2c5efede7b21f,64'h99bbdffb0e87c90e,64'h4c0d5f0a53516693,64'h9ed9501c02ff66bb,
64'hfe864c0d294cf1f4,64'h84b692405cc38f75,64'h3ba63dfd02b50fb8,64'h3e6ad357b0b7b45d,
64'h5a8dc374009ec4ed,64'h2b83b7ed95bb0790,64'h4c40695e0c29c9f3,64'he4f14ee68e6beb5c,
64'hc802df7a06ab5f9c,64'h141f2d137fd7081a,64'hc44812c9a6c91783,64'h28d6d652f210fc59,
64'h2eaeab70dee055c4,64'h9c7b4d0680d372ea,64'h7e7f303950029c3a,64'h5466ab558f6817fc,
64'hfc399005b810a2ef,64'h67cab0a01e964566,64'h86ac38ebe613b147,64'hfffffffec0000001,
64'h6a735604f3366569,64'h6dc5ae0d223eab16,64'ha11474afc1c4737f,64'hd0da26a62ace2fcf,
64'h98457f92844ad082,64'h9365f17424125b7a,64'hfcd96a63a536a724,64'h7522ed09dc17347b,
64'hfdc120f111d1e8f7,64'ha308326eabbc2cb5,64'h11b1ccfb83a19c03,64'hb8b13869db3a0094,
64'h4fb287f08e702149,64'ha0ab7e95c458c04e,64'h2df4571d7b3b7c4f,64'h57f14e8e202dad89,
64'h4a9a7006f9b48b31,64'h73519444cc5b0189,64'hb2dc621f68c63bd8,64'he11dff7751eaabb1,
64'hcc243b3d6da23b37,64'hb0dd08ecfbf7bc6c,64'hffab1c435b267edc,64'hef785c402fd58aba,
64'hdbd20d332b4b5e74,64'hf31566a7f1f722b4,64'hf2336dec512c82f9,64'h048d0b3a0d644547,
64'h027ba8f431f25136,64'h7d6fc1280e5c7125,64'h49d121a37e671e55,64'h0010000000000010,
64'h4c41efb63b6bc159,64'h0c46c44e398528a3,64'h4504295d6a2e396d,64'h09cd0976225e993f,
64'h2decfc45bb920c3f,64'ha769004743919df4,64'hb48144bbb33ad472,64'hc338d01992d4e785,
64'h37f658bdddbcf644,64'h53377bff21d0f922,64'ha981abe0aa6a2cd3,64'hb3db2a02e05fecd8,
64'h9fd0c98125299e3f,64'h7096d247ab9871ef,64'h0774c7bfa056a1f7,64'h67cd5a6a9616f68c,
64'h6b51b86e2013d89e,64'h057076fdb2b760f2,64'ha9880d2b2185393f,64'h9c9e29dc51cd7d6c,
64'h99005beec0d56bf4,64'hc283e5a1affae104,64'hb889025894d922f1,64'he51adac97e421f8c,
64'h85d5d56d9bdc0ab9,64'hd38f69a0101a6e5e,64'hcfcfe6066a005388,64'h8a8cd56a31ed0300,
64'h3f8732009702145e,64'h4cf95613c3d2c8ad,64'h30d5871d5cc27629,64'hfffffffef8000001,
64'hed4e6abfbe66ccae,64'h4db8b5c16447d563,64'h34228e95d8388e70,64'h3a1b44d4a559c5fa,
64'hd308aff190895a11,64'hd26cbe2dc4824b70,64'h9f9b2d4bf4a6d4e5,64'haea45da09b82e690,
64'h3fb8241e023a3d1f,64'h7461064d75778597,64'ha236399ed0743381,64'h9716270cbb674013,
64'he9f650fd31ce042a,64'h54156fd2788b180a,64'h25be8ae38f676f8a,64'heafe29d0e405b5b2,
64'he9534dffff369167,64'hee6a3287b98b6032,64'h165b8c43ed18c77b,64'hfc23bfee0a3d5577,
64'h398487678db44767,64'h961ba11d1f7ef78e,64'h9ff56387eb64cfdc,64'hddef0b8745fab158,
64'h9b7a41a5e5696bcf,64'h9e62acd47e3ee457,64'hfe466dbcaa259060,64'h2091a16721ac88a9,
64'h404f751e463e4a27,64'h6fadf824a1cb8e25,64'h693a24340fcce3cb,64'h0002000000000002,
64'he9883df5e76d782c,64'ha188d8892730a515,64'h68a0852b4d45c72e,64'h2139a12ea44bd328,
64'h25bd9f8897724188,64'h94ed2008687233bf,64'hd6902896b6675a8f,64'h78671a02d25a9cf1,
64'h86fecb173bb79ec9,64'hca66ef7f243a1f25,64'hb530357b754d459b,64'h167b65405c0bfd9b,
64'h33fa193004a533c8,64'h2e12da48d5730e3e,64'h20ee98f7d40ad43f,64'h8cf9ab4cd2c2ded2,
64'h4d6a370d84027b14,64'hc0ae0edef656ec1f,64'h353101a54430a728,64'h9393c53b0a39afae,
64'h93200b7d581aad7f,64'h98507cb3b5ff5c21,64'hf711204a329b245f,64'h9ca35b58afc843f2,
64'hf0babaacd37b8158,64'h5a71ed33c2034dcc,64'h19f9fcc0cd400a71,64'h11519aad463da060,
64'h47f0e63fd2e0428c,64'h699f2ac2187a5916,64'he61ab0e2cb984ec6,64'hfffffffeff000001,
64'h5da9cd57b7ccd996,64'ha9b716b78c88faad,64'h068451d2bb0711ce,64'hc7436899d4ab38c0,
64'hfa6115fd52112b43,64'h1a4d97c5b890496e,64'h73f365a91e94da9d,64'h15d48bb413705cd2,
64'h27f70483a04747a4,64'h2e8c20c98eaef0b3,64'hf446c732fa0e8671,64'hb2e2c4e0f76ce803,
64'hdd3eca1ee639c086,64'hca82adf98f116302,64'hc4b7d15bb1ecedf2,64'hdd5fc5395c80b6b7,
64'h3d2a69bfdfe6d22d,64'hddcd465037316c07,64'ha2cb7187dda318f0,64'h3f8477fda147aaaf,
64'h273090ecd1b688ed,64'h52c3742363efdef2,64'h93feac707d6c99fc,64'h1bbde170e8bf562b,
64'h336f48349cad2d7a,64'h33cc559a6fc7dc8b,64'h1fc8cdb79544b20c,64'he412342c04359116,
64'h2809eea3a8c7c945,64'h6df5bf04343971c5,64'had274485e1f99c7a,64'hc0003fff40000001,
64'h9d3107be3cedaf06,64'h74311b10c4e614a3,64'h4d1410a529a8b8e6,64'h04273425d4897a65,
64'h04b7b3f112ee4831,64'h329da400ed0e4678,64'h3ad20512b6cceb52,64'hef0ce33f7a4b539f,
64'hf0dfd9620776f3da,64'h794cddef848743e5,64'hb6a606aecea9a8b4,64'ha2cf6ca76b817fb4,
64'h067f43260094a679,64'h45c25b48daae61c8,64'h241dd31eda815a88,64'hd19f3568da585bdb,
64'h89ad46e130804f63,64'h3815c1dbbecadd84,64'h06a62034a88614e5,64'h527278a7214735f6,
64'h3264016f8b0355b0,64'hf30a0f9596bfeb85,64'h3ee224092653648c,64'hd3946b6a55f9087f,
64'h1e1757559a6f702b,64'h8b4e3da5f84069ba,64'he33f3f9739a8014f,64'h022a3355a8c7b40c,
64'h88fe1cc77a5c0852,64'h4d33e558030f4b23,64'h5cc3561c197309d9,64'hfffffffeffe00001,
64'h4bb539aab6f99b33,64'h7536e2d691911f56,64'h40d08a3a1760e23a,64'h18e86d133a956718,
64'hbf4c22bf0a422569,64'h4349b2f87712092e,64'h6e7e6cb4c3d29b54,64'hc2ba9175c26e0b9b,
64'h84fee08ff408e8f5,64'ha5d1841891d5de17,64'hfe88d8e57f41d0cf,64'hb65c589b7eed9d01,
64'h5ba7d9439cc73811,64'hd95055be71e22c61,64'hd896fa2ab63d9dbf,64'h3babf8a70b9016d7,
64'h67a54d379bfcda46,64'h3bb9a8c9e6e62d81,64'h14596e30fbb4631e,64'h27f08eff9428f556,
64'h64e6121d3a36d11e,64'hca586e83ac7dfbdf,64'h927fd58d8fad9340,64'ha377bc2d7d17eac6,
64'hc66de905d395a5b0,64'ha6798ab2adf8fb92,64'h83f919b672a89642,64'h5c8246854086b223,
64'h65013dd41518f929,64'h6dbeb7e026872e39,64'hd5a4e88ffc3f3390,64'hf80007ff08000001,
64'h53a620f7879db5e1,64'hae862361789cc295,64'h49a282146535171d,64'h6084e6845a912f4d,
64'he096f67d425dc907,64'h0653b4801da1c8cf,64'hc75a40a196d99d6b,64'h3de19c67cf496a74,
64'hde1bfb2b80eede7c,64'h6f299bbd9090e87d,64'h96d4c0d559d53517,64'h9459ed946d702ff7,
64'he0cfe863e01294d0,64'h08b84b691b55cc39,64'h0483ba63db502b51,64'hba33e6ac7b4b0b7c,
64'hb135a8db861009ed,64'h8702b83af7d95bb1,64'h60d4c4063510c29d,64'h4a4e4f14a428e6bf,
64'h064c802df1606ab6,64'h7e6141f252d7fd71,64'h87dc4480a4ca6c92,64'h3a728d6d2abf2110,
64'ha3c2eaea134dee06,64'hd169c7b3ff080d38,64'h3c67e7f2c735002a,64'h8045466a3518f682,
64'hd11fc3982f4b810b,64'ha9a67caa6061e965,64'heb986ac2a32e613c,64'hfffffffefffc0001,
64'ha976a734b6df3367,64'h4ea6dc5a923223eb,64'hc81a114682ec1c48,64'h031d0da26752ace3,
64'hf7e98457014844ae,64'h4869365ecee24126,64'h8dcfcd96187a536b,64'hb857522e184dc174,
64'h709fdc119e811d1f,64'h34ba3082f23abbc3,64'h3fd11b1c8fe83a1a,64'hf6cb8b128fddb3a1,
64'heb74fb279398e703,64'hfb2a0ab6ee3c458d,64'h3b12df4536c7b3b8,64'h27757f14c17202db,
64'h4cf4a9a6b37f9b49,64'he77735185cdcc5b1,64'h428b2dc5df768c64,64'h44fe11dfb2851eab,
64'h4c9cc2436746da24,64'h394b0dd0558fbf7c,64'h124ffab1b1f5b268,64'h546ef7856fa2fd59,
64'h18cdbd20ba72b4b6,64'hd4cf315595bf1f73,64'hd07f23360e5512c9,64'hab9048d00810d645,
64'heca027b9a2a31f26,64'hedb7d6fb24d0e5c8,64'h1ab49d11ff87e672,64'hff0000ff01000001,
64'hea74c41e10f3b6bd,64'h75d0c46bcf139853,64'h693450422ca6a2e4,64'h6c109cd02b5225ea,
64'h3c12decf884bb921,64'h20ca768fe3b4391a,64'hb8eb481392db33ae,64'h87bc338c79e92d4f,
64'h9bc37f64f01ddbd0,64'h6de5337752121d10,64'h32da981a8b3aa6a3,64'h328b3db26dae05ff,
64'h1c19fd0c7c02529a,64'he117096c436ab988,64'he090774b9b6a056b,64'h97467cd50f696170,
64'h7626b51b10c2013e,64'hf0e057067efb2b77,64'h6c1a988066a21854,64'h2949c9e274851cd8,
64'h40c990057e2c0d57,64'hefcc283d6a5affaf,64'hd0fb888f54994d93,64'h074e51ada557e422,
64'h54785d5d0269bdc1,64'h1a2d38f67fe101a7,64'hc78cfcfd98e6a006,64'hd008a8cc86a31ed1,
64'hba23f87265e97022,64'h7534cf94ec0c3d2d,64'h9d730d57d465cc28,64'hfffffffeffff8001,
64'h352ed4e676dbe66d,64'ha9d4db8ab246447e,64'h19034228d05d8389,64'ha063a1b3acea559d,
64'h5efd308aa0290896,64'h490d26cb99dc4825,64'hb1b9f9b2230f4a6e,64'h970aea454309b82f,
64'h2e13fb8213d023a4,64'ha697460fbe475779,64'hc7fa2362d1fd0744,64'hfed9716171fbb675,
64'hbd6e9f6452731ce1,64'h7f6541567dc788b2,64'h07625be8a6d8f677,64'ha4eeafe1f82e405c,
64'he99e9533f66ff36a,64'hfceee6a22b9b98b7,64'h885165b83beed18d,64'ha89fc23b5650a3d6,
64'h89939847ece8db45,64'h872961b98ab1f7f0,64'h0249ff56363eb64d,64'hea8ddeefcdf45fac,
64'h4319b7a3d74e5697,64'hba99e62a12b7e3ef,64'hfa0fe465e1caa25a,64'h75720919a1021ac9,
64'h5d9404f6f45463e5,64'h1db6fadf649a1cb9,64'hc35693a17ff0fccf,64'hffe0001f00200001,
64'h7d4e9883621e76d8,64'haeba188cd9e2730b,64'h8d268a07c594d45d,64'hcd821399456a44be,
64'he7825bd911097725,64'hc4194ed13c768724,64'h571d6902325b6676,64'h30f786716f3d25aa,
64'h13786fec9e03bb7a,64'h0dbca66eea4243a2,64'ha65b5302b16754d5,64'h265167b62db5c0c0,
64'hc3833fa0cf804a54,64'h1c22e12d886d5731,64'hbc120ee8d36d40ae,64'h12e8cf9aa1ed2c2e,
64'h4ec4d6a322184028,64'h3e1c0ae0afdf656f,64'h8d83530f8cd4430b,64'h0529393c4e90a39b,
64'h281932008fc581ab,64'h3df985078d4b5ff6,64'hba1f71114a9329b3,64'hc0e9ca34f4aafc85,
64'hea8f0baac04d37b9,64'h2345a71eaffc2035,64'h58f19f9f731cd401,64'hfa011518b0d463db,
64'hd7447f0d8cbd2e05,64'h6ea699f23d8187a6,64'h13ae61aafa8cb985,64'hfffffffefffff001,
64'h66a5da9c6edb7cce,64'h553a9b711648c890,64'he32068443a0bb072,64'h740c7436159d4ab4,
64'h4bdfa61114052113,64'h6921a4d9133b8905,64'h56373f360461e94e,64'h32e15d4888613706,
64'h85c27f6fc27a0475,64'hf4d2e8c117c8eaf0,64'h98ff446bda3fa0e9,64'h7fdb2e2bce3f76cf,
64'hf7add3ebaa4e639d,64'hcfeca82a0fb8f117,64'h20ec4b7cf4db1ecf,64'h949dd5fbbf05c80c,
64'hdd33d2a5becdfe6e,64'h3f9ddcd425737317,64'h710a2cb6a77dda32,64'h5513f8472aca147b,
64'h713273089d9d1b69,64'h10e52c3731563efe,64'h60493fea66c7d6ca,64'h9d51bbdd79be8bf6,
64'h286336f45ae9cad3,64'h37533cc52256fc7e,64'hdf41fc8bfc39544c,64'heeae41225420435a,
64'h6bb2809e7e8a8c7d,64'he3b6df5b0c934398,64'h386ad2740ffe1f9a,64'hfffc000300040001,
64'h0fa9d3106c43cedb,64'hb5d74310fb3c4e62,64'h71a4d14098b29a8c,64'h59b04272e8ad4898,
64'h7cf04b7ac2212ee5,64'h988329d9a78ed0e5,64'h4ae3ad20064b6ccf,64'hc61ef0cd6de7a4b6,
64'hc26f0dfcd3c07770,64'hc1b794cd1d484875,64'h74cb6a5ff62cea9b,64'h04ca2cf6c5b6b818,
64'h987067f399f0094b,64'he3845c24d10daae7,64'h578241dcda6da816,64'h425d19f3143da586,
64'h09d89ad464430805,64'h27c3815bf5fbecae,64'hb1b06a61519a8862,64'ha0a52726e9d21474,
64'ha503263f71f8b036,64'h47bf30a0b1a96bff,64'hb743ee2189526537,64'h781d39463e955f91,
64'hfd51e1747809a6f8,64'h6468b4e375ff8407,64'heb1e33f30e639a81,64'hbf4022a2761a8c7c,
64'h7ae88fe15197a5c1,64'h4dd4d33e07b030f5,64'h6275cc34ff519731,64'hfffffffefffffe01,
64'h4cd4bb534ddb6f9a,64'h0aa7536e22c91912,64'hdc640d07c741760f,64'h8e818e8642b3a957,
64'ha97bf4c18280a423,64'h6d24349ac2677121,64'h4ac6e7e6808c3d2a,64'h465c2ba8d10c26e1,
64'h70b84fed984f408f,64'h1e9a5d1822f91d5e,64'hf31fe88c9b47f41e,64'h2ffb65c559c7eeda,
64'h7ef5ba7d1549cc74,64'h39fd950521f71e23,64'h241d896f7e9b63da,64'h9293babef7e0b902,
64'h5ba67a5477d9bfce,64'h27f3bb9a64ae6e63,64'hce21459614efbb47,64'haaa27f0845594290,
64'hee264e6033b3a36e,64'h421ca586a62ac7e0,64'hcc0927fc8cd8fada,64'h53aa377b6f37d17f,
64'ha50c66ddeb5d395b,64'h46ea6798644adf90,64'h9be83f90ff872a8a,64'hddd5c8238a84086c,
64'h6d7650136fd15190,64'h1c76dbeb61926873,64'hc70d5a4dc1ffc3f4,64'hffff7fff80008001,
64'ha1f53a616d8879dc,64'hd6bae8615f6789cd,64'h8e349a2793165352,64'h0b36084e5d15a913,
64'h6f9e096ef84425dd,64'h7310653ad4f1da1d,64'h295c75a3e0c96d9a,64'h58c3de196dbcf497,
64'h184de1bf9a780eee,64'h7836f29943a9090f,64'hae996d4b5ec59d54,64'h0099459ed8b6d703,
64'hb30e0cfdd33e012a,64'h3c708b847a21b55d,64'h4af0483b5b4db503,64'h484ba33e2287b4b1,
64'h613b135a2c886101,64'h44f8702b3ebf7d96,64'hd6360d4b6a33510d,64'h9414a4e45d3a428f,
64'h54a064c7ae3f1607,64'h28f7e613f6352d80,64'h36e87dc4112a4ca7,64'hef03a727e7d2abf3,
64'h1faa3c2e8f0134df,64'h2c8d169c4ebff081,64'hfd63c67d81cc7351,64'h97e80453cec35190,
64'hef5d11fb4a32f4b9,64'h69ba9a6760f6061f,64'hec4eb985bfea32e7,64'hfffffffeffffffc1,
64'hc99a9769a9bb6df4,64'hc154ea6d04592323,64'h3b8c81a0d8e82ec2,64'h31d031d0a856752b,
64'hb52f7e9790501485,64'heda48692784cee25,64'hc958dcfc101187a6,64'he8cb85743a2184dd,
64'h2e1709fd9309e812,64'h43d34ba2c45f23ac,64'h5e63fd115368fe84,64'hc5ff6cb7eb38fddc,
64'h8fdeb74f22a9398f,64'ha73fb2a0043ee3c5,64'hc483b12d2fd36c7c,64'hd25277571efc1721,
64'h4b74cf4a4efb37fa,64'ha4fe7772ac95cdcd,64'h39c428b2a29df769,64'h15544fe108ab2852,
64'h5dc4c9cbc676746e,64'h084394b0d4c558fc,64'hd98124fed19b1f5c,64'h2a7546ef4de6fa30,
64'hb4a18cdb1d6ba72c,64'h08dd4cf30c895bf2,64'hd37d07f15ff0e552,64'h9bbab903f150810e,
64'h0daeca026dfa2a32,64'ha38edb7ccc324d0f,64'h98e1ab49383ff87f,64'hffffefff10001001,
64'h943ea74badb10f3c,64'h7ad75d0bcbecf13a,64'hd1c693443262ca6b,64'ha166c1092ba2b523,
64'h6df3c12d7f0884bc,64'h6e620ca6fa9e3b44,64'hc52b8eb3bc192db4,64'h2b187bc30db79e93,
64'h4309bc37b34f01de,64'h2f06de5308752122,64'h95d32da8ebd8b3ab,64'ha01328b33b16dae1,
64'hd661c19efa67c026,64'h678e11702f4436ac,64'ha95e0906cb69b6a1,64'he9097466e450f697,
64'hec27626a65910c21,64'h489f0e0527d7efb3,64'h7ac6c1a90d466a22,64'h3282949c6ba74852,
64'h2a940c98d5c7e2c1,64'h051efcc27ec6a5b0,64'h26dd0fb862254995,64'hbde074e45cfa557f,
64'h23f54785b1e0269c,64'he591a2d2a9d7fe11,64'hffac78ced0398e6b,64'h12fd008a79d86a32,
64'hfdeba23e89465e98,64'h2d37534ccc1ec0c4,64'h3d89d73097fd465d,64'hfffffffefffffff9,
64'h993352ecb5376dbf,64'hb82a9d4d008b2465,64'hc77190335b1d05d9,64'ha63a0639750acea6,
64'h76a5efd2920a0291,64'h7db490d1ef099dc5,64'h592b1b9f420230f5,64'h7d1970ae2744309c,
64'hc5c2e13ef2613d03,64'h887a6973d88be476,64'h8bcc7fa1aa6d1fd1,64'h98bfed967d671fbc,
64'h31fbd6e9c4552732,64'h74e7f653a087dc79,64'h9890762525fa6d90,64'hfa4a4eea03df82e5,
64'hc96e99e889df6700,64'h749fceedf592b9ba,64'he73885157453beee,64'hc2aa89fb6115650b,
64'h4bb8993938cece8e,64'h810872959a98ab20,64'h9b30249f5a3363ec,64'h054ea8dde9bcdf46,
64'h9694319ae3ad74e6,64'hc11ba99da1912b7f,64'hda6fa0fd6bfe1cab,64'h537757203e2a1022,
64'hc1b5d93f8dbf4547,64'h3471db6f798649a2,64'h331c35690707ff10,64'hfffffdff02000201,
64'h9287d4e8f5b621e8,64'hcf5aeba0b97d9e28,64'hba38d267e64c594e,64'hb42cd820857456a5,
64'h8dbe78252fe11098,64'h8dcc41945f53c769,64'h98a571d5f78325b7,64'ha5630f77c1b6f3d3,
64'h48613786b669e03c,64'hc5e0dbc9a10ea425,64'hb2ba65b47d7b1676,64'hf40265158762db5d,
64'h5acc38339f4cf805,64'h8cf1c22d85e886d6,64'hf52bc11ff96d36d5,64'h3d212e8cbc8a1ed3,
64'hfd84ec4c6cb22185,64'ha913e1c004fafdf7,64'hcf58d83461a8cd45,64'hc6505292cd74e90b,
64'he55281923ab8fc59,64'h00a3df984fd8d4b6,64'h64dba1f6ac44a933,64'h37bc0e9c6b9f4ab0,
64'h847ea8f0363c04d4,64'hfcb23459753affc3,64'hbff58f193a0731ce,64'hc25fa0108f3b0d47,
64'h1fbd7447d128cbd3,64'h85a6ea691983d819,64'h67b13ae5b2ffa8cc,64'hffffffff00000000,
64'h33266a5d76a6edb8,64'h770553a94011648d,64'hf8ee32058b63a0bc,64'h54c740c6eea159d5,
64'heed4bdf972414053,64'h6fb69219dde133b9,64'h6b2563738840461f,64'h8fa32e1544e88614,
64'hb8b85c273e4c27a1,64'h510f4d2e3b117c8f,64'hf1798ff3554da3fb,64'h9317fdb24face3f8,
64'hc63f7adc788aa4e7,64'hee9cfec99410fb90,64'h13120ec4a4bf4db2,64'h7f4949dce07bf05d,
64'h192dd33d113bece0,64'hce93f9dcfeb25738,64'h5ce710a26e8a77de,64'hb855513ecc22aca2,
64'h49771326e719d9d2,64'h10210e52b3531564,64'h936604936b466c7e,64'h40a9d51b7d379be9,
64'h52d286331c75ae9d,64'h3823753394322570,64'hbb4df41f0d7fc396,64'hca6eeae347c54205,
64'h3836bb27d1b7e8a9,64'hc68e3b6d2f30c935,64'h066386ad20e0ffe2,64'hffffffbf00400041,
64'h1250fa9d1eb6c43d,64'h19eb5d74172fb3c5,64'h57471a4cbcc98b2a,64'h76859b03b0ae8ad5,
64'h11b7cf04a5fc2213,64'hf1b98831abea78ee,64'h3314ae3a9ef064b7,64'hb4ac61ee5836de7b,
64'h890c26f056cd3c08,64'h78bc1b78d421d485,64'h56574cb64faf62cf,64'h7e804ca250ec5b6c,
64'h6b59870613e99f01,64'h519e384570bd10db,64'h7ea578239f2da6db,64'ha7a425d0f79143db,
64'h7fb09d892d964431,64'h35227c37e09f5fbf,64'h79eb1b062c3519a9,64'hb8ca0a51b9ae9d22,
64'hfcaa503167571f8c,64'h40147bf2c9fb1a97,64'hac9b743e35889527,64'h06f781d38d73e956,
64'h908fd51d86c7809b,64'hbf96468a8ea75ff9,64'h57feb1e2e740e63a,64'h384bf401f1e761a9,
64'ha3f7ae885a25197b,64'hf0b4dd4c43307b04,64'h8cf6275c365ff51a,64'h1fffffffe0000000,
64'h0664cd4baed4ddb7,64'h6ee0aa74c8022c92,64'h9f1dc640316c7418,64'h6a98e8187dd42b3b,
64'hbdda97be8e48280b,64'hedf6d2425bbc2678,64'h2d64ac6e510808c4,64'h91f465c2289d10c3,
64'hf7170b8407c984f5,64'h2a21e9a5a7622f92,64'hbe2f31fdcaa9b480,64'h1262ffb649f59c7f,
64'h38c7ef5b6f11549d,64'h1dd39fd932821f72,64'hc26241d7d497e9b7,64'h6fe9293b3c0f7e0c,
64'h0325ba67a2277d9c,64'h19d27f3b9fd64ae7,64'h4b9ce2140dd14efc,64'hd70aaa2719845595,
64'hc92ee2641ce33b3b,64'h820421c9d66a62ad,64'h526cc0922d68cd90,64'he8153aa28fa6f37e,
64'h6a5a50c6038eb5d4,64'h07046ea6728644ae,64'h5769be83a1aff873,64'h794ddd5c08f8a841,
64'he706d7641a36fd16,64'h78d1c76d45e61927,64'hc0cc70d4e41c1ffd,64'hfffffff700080009,
64'h624a1f5343d6d888,64'h633d6bae22e5f679,64'hcae8e348d7993166,64'h6ed0b3601615d15b,
64'ha236f9dff4bf8443,64'h5e373105f57d4f1e,64'h266295c733de0c97,64'hb6958c3d2b06dbd0,
64'h112184de0ad9a781,64'h6f17836eba843a91,64'h2acae996a9f5ec5a,64'h8fd00993ca1d8b6e,
64'hed6b30dfe27d33e1,64'haa33c7080e17a21c,64'hafd4af03d3e5b4dc,64'hb4f484b97ef2287c,
64'heff613b045b2c887,64'h26a44f86dc13ebf8,64'hef3d635fe586a336,64'hd71941497735d3a5,
64'h9f954a05aceae3f2,64'h28028f7e393f6353,64'h35936e87a6b112a5,64'h40def03a31ae7d2b,
64'hb211faa310d8f014,64'hf7f2c8d071d4ec00,64'hcaffd63b9ce81cc8,64'he7097e7f5e3cec36,
64'hb47ef5d06b44a330,64'h9e169ba908660f61,64'hd19ec4eac6cbfea4,64'h03fffffffc000000,
64'h20cc99a955da9bb7,64'hcddc154dd9004593,64'h13e3b8c8062d8e83,64'had531d026fba8568,
64'hb7bb52f731c90502,64'h1dbeda484b7784cf,64'h85ac958d4a210119,64'hb23e8cb7a513a219,
64'h7ee2e17020f9309f,64'hc5443d33f4ec45f3,64'h17c5e63fb9553690,64'h224c5ff6a93eb390,
64'h6718fdeb0de22a94,64'hc3ba73fa665043ef,64'h384c483ada92fd37,64'h8dfd2526e781efc2,
64'h8064b74c7444efb4,64'h233a4fe753fac95d,64'h89739c4201ba29e0,64'h7ae1554483308ab3,
64'hb925dc4be39c6768,64'h70408438dacd4c56,64'h0a4d981245ad19b2,64'h5d02a75411f4de70,
64'h8d4b4a184071d6bb,64'h40e08dd48e50c896,64'haaed37cfd435ff0f,64'hef29bbaaa11f1509,
64'h5ce0daec4346dfa3,64'h2f1a38ed88bcc325,64'h78198e1a3c838400,64'hfffffffe00010002,
64'h0c4943ea687adb11,64'hec67ad74e45cbed0,64'h595d1c68daf3262d,64'hadda166b62c2ba2c,
64'hb446df3b5e97f089,64'h4bc6e6207eafa9e4,64'h24cc52b8c67bc193,64'h16d2b187a560db7a,
64'he224309ae15b34f1,64'hede2f06cf7508753,64'hc5595d32153ebd8c,64'h51fa01323943b16e,
64'hfdad661b1c4fa67d,64'h954678e081c2f444,64'h95fa95dffa7cb69c,64'h969e9096afde4510,
64'h3dfec275e8b65911,64'h04d489f0db827d7f,64'h5de7ac6bbcb0d467,64'h7ae32828cee6ba75,
64'hd3f2a93ff59d5c7f,64'ha50051ef2727ec6b,64'h66b26dd094d62255,64'ha81bde06a635cfa6,
64'h96423f53e21b1e03,64'h1efe591a0e3a9d80,64'h195ffac7739d0399,64'h5ce12fcfabc79d87,
64'h168fdeba0d689466,64'hf3c2d374410cc1ed,64'h9a33d89cd8d97fd5,64'h007fffffff800000,
64'h241993350abb5377,64'hb9bb82a91b2008b3,64'ha27c771860c5b1d1,64'h15aa63a04df750ad,
64'hd6f76a5e263920a1,64'h23b7db48e96ef09a,64'hf0b592b0c9442024,64'hf647d19614a27444,
64'h2fdc5c2de41f2614,64'hb8a887a5de9d88bf,64'h02f8bcc7f72aa6d2,64'h04498bfed527d672,
64'h8ce31fbce1bc4553,64'h38774e7f2cca087e,64'h270989073b525fa7,64'hd1bfa4a41cf03df9,
64'h900c96e90e889df7,64'h646749fc8a7f592c,64'h112e73884037453c,64'haf5c2aa7f0661157,
64'h1724bb897c738ced,64'h4e081086db59a98b,64'hc149b30188b5a337,64'h0ba054ea823e9bce,
64'hb1a96942680e3ad8,64'h481c11ba51ca1913,64'h355da6f9da86bfe2,64'hfde537747423e2a2,
64'hab9c1b5ce868dbf5,64'h65e3471d51179865,64'h0f0331c347907080,64'hdfffffff00002001,
64'he189287c6d0f5b63,64'h1d8cf5ae9c8b97da,64'h6b2ba38cbb5e64c6,64'h95bb42ccec585746,
64'hf688dbe68bd2fe12,64'h8978dcc38fd5f53d,64'ha4998a5678cf7833,64'hc2da563034ac1b70,
64'hfc4486127c2b669f,64'hbdbc5e0cfeea10eb,64'h98ab2ba5c2a7d7b2,64'h4a3f40260728762e,
64'h7fb5acc30389f4d0,64'h92a8cf1b90385e89,64'h92bf52bb7f4f96d4,64'h12d3d212d5fbc8a2,
64'he7bfd84ddd16cb23,64'h209a913dfb704fb0,64'h2bbcf58d57961a8d,64'h6f5c6504b9dcd74f,
64'h3a7e5527deb3ab90,64'hb4a00a3d44e4fd8e,64'h6cd64db9b29ac44b,64'h55037bc094c6b9f5,
64'hb2c847e9dc4363c1,64'h03dfcb2341c753b0,64'he32bff580e73a074,64'h2b9c25f9d578f3b1,
64'h42d1fbd701ad128d,64'h7e785a6e2821983e,64'h73467b133b1b2ffb,64'h000ffffffff00000,
64'h2483326681576a6f,64'hb737705483640117,64'hf44f8ee22c18b63b,64'h62b54c73a9beea16,
64'hfadeed4ae4c72415,64'hc476fb685d2dde14,64'h9e16b25599288405,64'h9ec8fa3242944e89,
64'h85fb8b853c83e4c3,64'h371510f49bd3b118,64'hc05f17983ee554db,64'hc089317f1aa4facf,
64'hb19c63f6fc3788ab,64'h470ee9cfa5994110,64'h24e13120c76a4bf5,64'hfa37f493a39e07c0,
64'h320192dd01d113bf,64'h8c8ce93f114feb26,64'h8225ce708806e8a8,64'h35eb8554de0cc22b,
64'h62e49770cf8e719e,64'ha9c102103b6b3532,64'h382936601116b467,64'h41740a9d1047d37a,
64'h16352d284d01c75b,64'ha9038236aa394323,64'hc6abb4de7b50d7fd,64'hdfbca6edce847c55,
64'h7573836b3d0d1b7f,64'h6cbc68e34a22f30d,64'h01e0663868f20e10,64'hfbffffff00000401,
64'hbc31250eeda1eb6d,64'hc3b19eb5139172fc,64'h4d657471576bcc99,64'h52b768595d8b0ae9,
64'hded11b7c117a5fc3,64'h712f1b9811fabea8,64'hb493314a2f19ef07,64'h185b4ac60695836e,
64'h3f8890c22f856cd4,64'hb7b78bc0ffdd421e,64'hd3156573f854faf7,64'h4947e80480e50ec6,
64'h0ff6b59860713e9a,64'hf25519e292070bd2,64'h9257ea56efe9f2db,64'hc25a7a419abf7915,
64'hbcf7fb091ba2d965,64'h04135227bf6e09f6,64'h65779eb14af2c352,64'h2deb8ca0773b9aea,
64'h074fcaa4fbd67572,64'h56940147689c9fb2,64'had9ac9b69653588a,64'h6aa06f77b298d73f,
64'hf65908fc5b886c79,64'h007bf9646838ea76,64'h9c657fea81ce740f,64'he57384be5aaf1e77,
64'h685a3f7a8035a252,64'h4fcf0b4d85043308,64'hae68cf61c7636600,64'h0001fffffffe0000,
64'h2490664cb02aed4e,64'h36e6ee0a706c8023,64'hbe89f1dba58316c8,64'h4c56a98e3537dd43,
64'h7f5bdda8fc98e483,64'h988edf6c8ba5bbc3,64'h73c2d64a53251081,64'hf3d91f45685289d2,
64'hb0bf717007907c99,64'h06e2a21e937a7623,64'hb80be2f267dcaa9c,64'h3811262fc3549f5a,
64'hb6338c7e3f86f116,64'h08e1dd39f4b32822,64'h649c2623b8ed497f,64'h1f46fe927473c0f8,
64'h2640325b803a2278,64'h51919d27a229fd65,64'h1044b9ce1100dd15,64'ha6bd70a9fbc19846,
64'h4c5c92edd9f1ce34,64'hd5382041476d66a7,64'h270526cbe222d68d,64'hc82e8152e208fa70,
64'ha2c6a5a469a038ec,64'hb520704635472865,64'h78d5769b6f6a1b00,64'h7bf794dd59d08f8b,
64'h2eae706d47a1a370,64'h6d978d1c09445e62,64'h003c0cc70d1e41c2,64'hff7fffff00000081,
64'h778624a17db43d6e,64'h987633d622722e60,64'he9acae8d4aed7994,64'hea56ed0a4bb1615e,
64'hbbda236ee22f4bf9,64'h0e25e373023f57d5,64'h3692662925e33de1,64'h430b695880d2b06e,
64'h87f11217c5f0ad9b,64'h56f6f177dffba844,64'h3a62acae5f0a9f5f,64'h4928fd00501ca1d9,
64'hc1fed6b24c0e27d4,64'hde4aa33b9240e17b,64'hb24afd4a3dfd3e5c,64'h784b4f47d357ef23,
64'h779eff60c3745b2d,64'h40826a44b7edc13f,64'hccaef3d5695e586b,64'hc5bd71934ee7735e,
64'hc0e9f953df7aceaf,64'hcad280282d1393f7,64'hd5b3593612ca6b12,64'h2d540deed6531ae8,
64'hfecb211eab710d90,64'h400f7f2c4d071d4f,64'h338caffd3039ce82,64'h3cae7097ab55e3cf,
64'hcd0b47ee9006b44b,64'h09f9e169b0a08661,64'h15cd19ec38ec6cc0,64'h00003fffffffc000,
64'h44920cc956055daa,64'ha6dcddc0ae0d9005,64'h17d13e3b74b062d9,64'ha98ad53126a6fba9,
64'hafeb7bb47f931c91,64'hb311dbecf174b779,64'hee785ac86a64a211,64'hde7b23e7ed0a513b,
64'hf617ee2d20f20f94,64'ha0dc5443326f4ec5,64'h97017c5dccfb9554,64'hc70224c5386a93ec,
64'h56c6718f87f0de23,64'hc11c3ba67e966505,64'h2c9384c4571da930,64'h03e8dfd24e8e781f,
64'h04c8064b7007444f,64'h6a3233a494453fad,64'h6208973962201ba3,64'h54d7ae14ff783309,
64'h898b925d3b3e39c7,64'h3aa7040808edacd5,64'h64e0a4d91c445ad2,64'h1905d02a5c411f4e,
64'h9458d4b40d34071e,64'h76a40e0866a8e50d,64'h0f1aaed36ded4360,64'haf7ef29b0b3a11f2,
64'h05d5ce0da8f4346e,64'hcdb2f1a2c1288bcd,64'hc007819821a3c839,64'hffefffff00000011,
64'h4ef0c493efb687ae,64'h130ec67ac44e45cc,64'h9d3595d1295daf33,64'h5d4adda109762c2c,
64'hf77b446cfc45e980,64'h61c4bc6e0047eafb,64'he6d24cc444bc67bd,64'h48616d2ad01a560e,
64'hb0fe224258be15b4,64'h8adede2e7bff7509,64'h274c5595abe153ec,64'he9251f9f2a03943c,
64'h983fdad5c981c4fb,64'hbbc95466d2481c30,64'h96495fa8c7bfa7cc,64'haf0969e85a6afde5,
64'h6ef3dfebb86e8b66,64'h28104d4876fdb828,64'hb995de7a0d2bcb0e,64'h58b7ae3229dcee6c,
64'h381d3f2a5bef59d6,64'h395a5004e5a2727f,64'hdab66b2602594d63,64'h05aa81bddaca635d,
64'h1fd96423d56e21b2,64'h2801efe569a0e3aa,64'hc67195fee60739d1,64'h2795ce12d56abc7a,
64'hb9a168fd3200d68a,64'he13f3c2c561410cd,64'h02b9a33d871d8d98,64'h000007fffffff800,
64'hc89241986ac0abb6,64'h74db9bb7b5c1b201,64'he2fa27c68e960c5c,64'hf5315aa544d4df76,
64'hf5fd6f75aff26393,64'hf6623b7cbe2e96f0,64'hfdcf0b582d4c9443,64'hbbcf647c5da14a28,
64'h9ec2fdc5241e41f3,64'h741b8a88064de9d9,64'h92e02f8b399f72ab,64'h98e04498270d527e,
64'haad8ce3150fe1bc5,64'h782387746fd2cca1,64'h059270988ae3b526,64'h207d1bfa29d1cf04,
64'h209900c94e00e88a,64'h6d4646743288a7f6,64'hac4112e68c440375,64'hea9af5c1bfef0662,
64'h3131724b8767c739,64'h6754e080a11db59b,64'hcc9c149a63888b5b,64'h4320ba050b8823ea,
64'h528b1a9641a680e4,64'h6ed481c0acd51ca2,64'h01e355da6dbda86c,64'hd5efde52a167423f,
64'h40bab9c1751e868e,64'h79b65e33f825117a,64'hf800f03224347908,64'hfffdffff00000003,
64'h49de18923df6d0f6,64'h8261d8ced889c8ba,64'hb3a6b2b9852bb5e7,64'h8ba95bb3a12ec586,
64'h1eef688d9f88bd30,64'hac38978d2008fd60,64'h7cda499828978cf8,64'h490c2da51a034ac2,
64'h961fc447cb17c2b7,64'hf15bdbc4ef7feea2,64'h84e98ab2357c2a7e,64'h9d24a3f365407288,
64'hb307fb5a193038a0,64'h17792a8cda490386,64'h92c92bf498f7f4fa,64'h75e12d3cab4d5fbd,
64'h4dde7bfd370dd16d,64'h050209a90edfb705,64'h5732bbcf01a57962,64'h8b16f5c5c53b9dce,
64'h4703a7e50b7deb3b,64'h272b4a007cb44e50,64'hbb56cd64204b29ad,64'h60b550375b594c6c,
64'hc3fb2c83baadc437,64'hc5003dfbed341c76,64'hf8ce32befcc0e73b,64'hc4f2b9c19aad5790,
64'hd7342d1ee6401ad2,64'h7c27e7852ac2821a,64'h00573467b0e3b1b3,64'h000000ffffffff00,
64'h59124832cd581577,64'hee9b737616b83641,64'h9c5f44f851d2c18c,64'h5ea62b54689a9bef,
64'hbebfadee15fe4c73,64'h1ecc476f97c5d2de,64'hbfb9e16a65a99289,64'h1779ec8f8bb42945,
64'hb3d85fb80483c83f,64'hee83715020c9bd3c,64'hb25c05f0c733ee56,64'h531c0892c4e1aa50,
64'h755b19c5ca1fc379,64'hef0470edadfa5995,64'h40b24e12d15c76a5,64'h840fa37ec53a39e1,
64'hc413201869c01d12,64'h4da8c8ce465114ff,64'h7588225c7188806f,64'hdd535eb777fde0cd,
64'he6262e4890ecf8e8,64'hacea9c0f7423b6b4,64'hb9938292ac71116c,64'hc864173fe171047e,
64'h8a5163524834d01d,64'hcdda9037559aa395,64'h803c6abacdb7b50e,64'h3abdfbca342ce848,
64'h48175737eea3d0d2,64'hcf36cbc5bf04a230,64'h1f001e0644868f21,64'hbfffbfff40000001,
64'h493bc31207beda1f,64'hd04c3b191b113918,64'h3674d65710a576bd,64'h51752b763425d8b1,
64'h03dded11b3f117a6,64'h158712f1a4011fac,64'h0f9b49330512f19f,64'hc92185b3e3406959,
64'h32c3f888d962f857,64'hde2b7b77ddeffdd5,64'h509d315606af8550,64'h13a4947e6ca80e51,
64'h1660ff6b43260714,64'h42ef25515b492071,64'hd259257dd31efea0,64'h6ebc25a73569abf8,
64'h69bbcf7f46e1ba2e,64'h60a04134c1dbf6e1,64'hcae657792034af2d,64'h5162deb878a773ba,
64'ha8e074fc016fbd68,64'h04e569400f9689ca,64'h776ad9ac24096536,64'h8c16aa066b6b298e,
64'h387f65905755b887,64'h58a007bf3da6838f,64'hbf19c6573f981ce8,64'h189e57383355aaf2,
64'hdae685a31cc8035b,64'hcf84fcefe5585044,64'ha00ae68c561c7637,64'h0000001fffffffe0,
64'h2b22490639ab02af,64'hfdd36e6de2d706c9,64'h938be89e8a3a5832,64'h2bd4c56a6d13537e,
64'hb7d7f5bd22bfc98f,64'h43d988edb2f8ba5c,64'hf7f73c2c6cb53252,64'h62ef3d9191768529,
64'h367b0bf6e0907908,64'h9dd06e29841937a8,64'h564b80bdd8e67dcb,64'h0a638112589c354a,
64'heeab6337d943f870,64'h7de08e1d55bf4b33,64'h681649c1fa2b8ed5,64'hf081f46ef8a7473d,
64'hd88264024d3803a3,64'h29b51919a8ca22a0,64'h2eb1044b6e31100e,64'h7baa6bd68effbc1a,
64'h1cc4c5c9121d9f1d,64'h959d53816e8476d7,64'h97327051d58e222e,64'h590c82e7bc2e2090,
64'h714a2c69e9069a04,64'h79bb52068ab35473,64'h50078d5719b6f6a2,64'h0757bf7946859d09,
64'hc902eae63dd47a1b,64'h19e6d978b7e09446,64'he3e003bfe890d1e5,64'hf7fff7ff08000001,
64'h2927786220f7db44,64'h1a09876323622723,64'h66ce9aca8214aed8,64'hea2ea56de684bb17,
64'h407bbda1f67e22f5,64'h82b0e25db48023f6,64'h21f3692640a25e34,64'hf92430b59c680d2c,
64'h26587f10fb2c5f0b,64'h7bc56f6e9bbdffbb,64'h0a13a62ac0d5f0aa,64'he274928eed9501cb,
64'h82cc1fece864c0e3,64'he85de4a94b69240f,64'h1a4b24afba63dfd4,64'h0dd784b4e6ad357f,
64'h4d3779efa8dc3746,64'hec140825b83b7edd,64'h795ccaeec40695e6,64'hca2c5bd64f14ee78,
64'h151c0e9f802df7ad,64'hc09cad2741f2d13a,64'h4eed5b3544812ca7,64'h5182d5408d6d6532,
64'h270fecb1eaeab711,64'h2b1400f7c7b4d072,64'h17e338cae7f3039d,64'hc313cae6466ab55f,
64'hbb5cd0b3c399006c,64'h99f09f9d7cab0a09,64'h34015cd16ac38ec7,64'h00000003fffffffc,
64'h25644920a7356056,64'hffba6dccdc5ae0da,64'hd2717d1311474b07,64'h457a98ad0da26a70,
64'h36fafeb78457f932,64'h887b311d365f174c,64'hdefee784cd96a64b,64'hec5de7b1522ed0a6,
64'h06cf617edc120f21,64'h13ba0dc5308326f5,64'haac970171b1ccfba,64'hc14c70218b1386aa,
64'h1dd56c66fb287f0e,64'hafbc11c30ab7e967,64'h6d02c937df4571db,64'h7e103e8d7f14e8e8,
64'hbb104c7fa9a70075,64'h0536a32335194454,64'h45d620892dc62202,64'hcf754d7a11dff784,
64'h639898b8c243b3e4,64'h32b3aa700dd08edb,64'h52e64e09fab1c446,64'h0b21905cf785c412,
64'h8e29458cbd20d341,64'haf376a4031566a8f,64'hca00f1aa2336ded5,64'he0eaf7ee48d0b3a2,
64'hb9205d5c27ba8f44,64'h433cdb2ed6fc1289,64'h7c7c00779d121a3d,64'hfefffeff01000001,
64'h8524ef0bc41efb69,64'ha34130ebc46c44e5,64'h0cd9d359504295db,64'h3d45d4ad9cd09763,
64'h680f77b3decfc45f,64'h50561c4b7690047f,64'h843e6d2448144bc7,64'h9f248616338d01a6,
64'ha4cb0fe17f658be2,64'haf78aded3377bff8,64'hc14274c4981abe16,64'hbc4e92513db2a03a,
64'hb05983fcfd0c981d,64'h3d0bbc95096d2482,64'h83496495774c7bfb,64'h21baf0967cd5a6b0,
64'h49a6ef3db51b86e9,64'h7d82810457076fdc,64'h4f2b995d9880d2bd,64'h19458b7ac9e29dcf,
64'h62a381d39005bef6,64'hd81395a4283e5a28,64'h29ddab6688902595,64'hca305aa751adaca7,
64'he4e1fd955d5d56e3,64'hc562801e38f69a0f,64'h62fc6718fcfe6074,64'h3862795ca8cd56ac,
64'h976b9a15f873200e,64'hf33e13f2cf956142,64'h26802b9a0d5871d9,64'h8000000000000000,
64'h44ac8923d4e6ac0b,64'hdff74db8db8b5c1c,64'h3a4e2fa24228e961,64'h08af5315a1b44d4e,
64'hc6df5fd6308aff27,64'h910f662326cbe2ea,64'hbbdfdceff9b2d4ca,64'h5d8bbcf5ea45da15,
64'he0d9ec2efb8241e5,64'h627741b8461064df,64'hd5592e02236399f8,64'hd8298e03716270d6,
64'h43baad8c9f650fe2,64'h35f782384156fd2d,64'hada059265be8ae3c,64'h0fc207d1afe29d1d,
64'h7762098f9534e00f,64'h80a6d463e6a3288b,64'hc8bac41065b8c441,64'h99eea9aec23bfef1,
64'h8c7313169848767d,64'ha656754d61ba11dc,64'h4a5cc9c0ff563889,64'hc164320adef0b883,
64'hf1c528b0b7a41a69,64'h35e6ed47e62acd52,64'h79401e34e466dbdb,64'hdc1d5efd091a1675,
64'h97240bab04f751e9,64'he8679b64fadf8252,64'h6f8f800e93a24348,64'hffdfffdf00200001,
64'hf0a49de09883df6e,64'h7468261d188d889d,64'ha19b3a6a8a0852bc,64'ha7a8ba95139a12ed,
64'h2d01eef65bd9f88c,64'h2a0ac3894ed20090,64'h3087cda469028979,64'h53e490c28671a035,
64'hd49961fb6fecb17d,64'h15ef15bda66ef7ff,64'h58284e98530357c3,64'hd789d24967b65408,
64'h760b307f3fa19304,64'hc7a17791e12da491,64'hb0692c920ee98f80,64'h04375e12cf9ab4d6,
64'he934dde6d6a370de,64'h8fb050200ae0edfc,64'h69e5732b53101a58,64'h2328b16f393c53ba,
64'h4c54703a3200b7df,64'h1b0272b48507cb45,64'h653bb56c711204b3,64'h39460b54ca35b595,
64'hbc9c3fb20babaadd,64'h38ac5003a71ed342,64'h8c5f8ce29f9fcc0f,64'h870c4f2b1519aad6,
64'h52ed73427f0e6402,64'hde67c27d99f2ac29,64'he4d0057261ab0e3c,64'h1000000000000000,
64'ha8959123da9cd582,64'h9bfee9b69b716b84,64'he749c5f368451d2d,64'h4115ea62743689aa,
64'h38dbebfaa6115fe5,64'hd221ecc3a4d97c5e,64'hd77bfb9d3f365a9a,64'h6bb1779e5d48bb43,
64'h7c1b3d857f70483d,64'h2c4ee836e8c20c9c,64'h1aab25c0446c733f,64'h5b0531c02e2c4e1b,
64'hc87755b0d3eca1fd,64'h66bef046a82adfa6,64'h95b40b244b7d15c8,64'h61f840f9d5fc53a4,
64'h2eec4131d2a69c02,64'hb014da8bdcd46512,64'hf91758812cb71889,64'hf33dd534f8477fdf,
64'h718e626273090ed0,64'h94cacea92c37423c,64'he94b99373feac712,64'hb82c8640bbde1711,
64'hfe38a51536f4834e,64'hc6bcdda83cc559ab,64'haf2803c5fc8cdb7c,64'h7b83abdf412342cf,
64'hf2e48174809eea3e,64'hdd0cf36bdf5bf04b,64'h0df1f001d2744869,64'hfffbfffb00040001,
64'h5e1493bbd3107bee,64'h6e8d04c34311b114,64'h9433674cd1410a58,64'h74f517524273425e,
64'h85a03dde4b7b3f12,64'h0541587129da4012,64'he610f9b3ad205130,64'h6a7c9217f0ce3407,
64'h7a932c3f0dfd9630,64'h22bde2b794cddf00,64'hab0509d26a606af9,64'h1af13a492cf6ca81,
64'h8ec1660f67f43261,64'hf8f42ef15c25b493,64'h160d259241dd31f0,64'h4086ebc219f3569b,
64'h5d269bbc9ad46e1c,64'h91f60a03815c1dc0,64'h0d3cae656a62034b,64'hc465162d27278a78,
64'h298a8e07264016fc,64'h63604e5630a0f969,64'haca776acee224097,64'h6728c16a3946b6b3,
64'h779387f5e175755c,64'hc71589ffb4e3da69,64'h318bf19c33f3f982,64'h50e189e522a3355b,
64'hca5dae678fe1cc81,64'hfbccf84ed33e5586,64'h9c9a00adcc3561c8,64'h0200000000000000,
64'hd512b223bb539ab1,64'h937fdd36536e2d71,64'h7ce938be0d08a3a6,64'hc822bd4b8e86d136,
64'h671b7d7ef4c22bfd,64'h5a443d98349b2f8c,64'hdaef7f72e7e6cb54,64'had762ef32ba91769,
64'h6f8367b04fee0908,64'h8589dd065d184194,64'h235564b7e88d8e68,64'hab60a63765c589c4,
64'h790eeab5ba7d9440,64'h4cd7de0895055bf5,64'h12b68164896fa2b9,64'h8c3f081ebabf8a75,
64'hc5dd88257a54d381,64'hd6029b50bb9a8ca3,64'hff22eb0f4596e312,64'h3e67baa67f08effc,
64'h0e31cc4c4e6121da,64'h929959d4a586e848,64'hdd29732627fd58e3,64'hf70590c7377bc2e3,
64'h5fc714a266de906a,64'hb8d79bb46798ab36,64'h95e500783f919b70,64'h2f70757bc824685a,
64'h5e5c902e5013dd48,64'hbba19e6cdbeb7e0a,64'he1be3dff5a4e890e,64'hffff7ffe80008001,
64'h4bc292773a620f7e,64'h8dd1a097e8623623,64'h12866ce99a28214b,64'h4e9ea2ea084e684c,
64'hd0b407bb096f67e3,64'hc0a82b0d653b4803,64'h1cc21f3675a40a26,64'h2d4f9242de19c681,
64'h0f526587e1bfb2c6,64'h0457bc56f299bbe0,64'hf560a1396d4c0d60,64'he35e2748459ed951,
64'hf1d82cc10cfe864d,64'hbf1e85dd8b84b693,64'h02c1a4b2483ba63e,64'ha810dd77a33e6ad4,
64'h8ba4d377135a8dc4,64'h123ec140702b83b8,64'ha1a795cc0d4c406a,64'h188ca2c5a4e4f14f,
64'h853151c064c802e0,64'hec6c09c9e6141f2e,64'h3594eed57dc44813,64'hace5182ca728d6d7,
64'h8ef270fe3c2eaeac,64'hf8e2b13f169c7b4e,64'hc6317e32c67e7f31,64'haa1c313c045466ac,
64'hf94bb5cc11fc3991,64'h5f799f099a67cab1,64'h13934015b986ac39,64'h0040000000000000,
64'hfaa25643976a7357,64'hf26ffba5ea6dc5af,64'h4f9d271781a11475,64'h590457a931d0da27,
64'h6ce36faf7e984580,64'h8b4887b2869365f2,64'h9b5defeddcfcd96b,64'hf5aec5dd857522ee,
64'h0df06cf609fdc121,64'h90b13ba04ba30833,64'h046aac96fd11b1cd,64'h956c14c66cb8b139,
64'h0f21dd56b74fb288,64'h699afbc0b2a0ab7f,64'he256d02bb12df458,64'h7187e1037757f14f,
64'hf8bbb103cf4a9a71,64'hbac0536977735195,64'hdfe45d6128b2dc63,64'h87ccf7544fe11e00,
64'hc1c63988c9cc243c,64'h12532b3a94b0dd09,64'hbba52e6424ffab1d,64'hbee0b21846ef785d,
64'hcbf8e2938cdbd20e,64'h571af3764cf31567,64'h12bca00f07f2336e,64'hc5ee0eaeb9048d0c,
64'h0bcb9205ca027ba9,64'hd77433ccdb7d6fc2,64'h5c37c7bfab49d122,64'hffffeffef0001001,
64'h4978524ea74c41f0,64'hb1ba34125d0c46c5,64'ha250cd9c9345042a,64'h89d3d45cc109cd0a,
64'hba1680f6c12decfd,64'hb81505610ca76901,64'h439843e68eb48145,64'he5a9f2477bc338d1,
64'h41ea4cb0bc37f659,64'h008af78ade53377c,64'h1eac14272da981ac,64'hfc6bc4e828b3db2b,
64'h7e3b0597c19fd0ca,64'hb7e3d0bb117096d3,64'h40583496090774c8,64'h95021bae7467cd5b,
64'h91749a6e626b51b9,64'h0247d8280e057077,64'hd434f2b8c1a9880e,64'h23119458949c9e2a,
64'h10a62a380c99005c,64'h5d8d8138fcc283e6,64'ha6b29dda0fb88903,64'h359ca30574e51adb,
64'h91de4e1f4785d5d6,64'h5f1c5627a2d38f6a,64'hf8c62fc578cfcfe7,64'h95438627008a8cd6,
64'hff2976b8a23f8733,64'hebef33e0534cf957,64'he2726801d730d588,64'h0008000000000000,
64'h3f544ac852ed4e6b,64'h3e4dff749d4db8b6,64'h69f3a4e29034228f,64'h2b208af5063a1b45,
64'h0d9c6df5efd308b0,64'hd16910f590d26cbf,64'hb36bbdfd1b9f9b2e,64'h5eb5d8bb70aea45e,
64'he1be0d9de13fb825,64'hb216277369746107,64'h608d55927fa2363a,64'hf2ad8297ed971628,
64'h01e43baad6e9f651,64'h2d335f77f6541570,64'h1c4ada057625be8b,64'h2e30fc204eeafe2a,
64'hff17761f99e9534f,64'h77580a6cceee6a33,64'hbbfc8bab85165b8d,64'h10f99eea89fc23c0,
64'h9838c73099398488,64'he24a656672961ba2,64'h7774a5cc249ff564,64'h77dc1642a8ddef0c,
64'h597f1c52319b7a42,64'h2ae35e6ea99e62ad,64'h42579401a0fe466e,64'h98bdc1d5572091a2,
64'he179723fd9404f76,64'hdaee8678db6fadf9,64'hcb86f8f735693a25,64'hfffffdfefe000201,
64'h092f0a49d4e9883e,64'h76374681eba188d9,64'hd44a19b2d268a086,64'hd13a7a8ad82139a2,
64'h7742d01e7825bda0,64'hf702a0ab4194ed21,64'h6873087c71d69029,64'hfcb53e480f78671b,
64'he83d49953786fecc,64'h80115ef0dbca66f0,64'h83d5828465b53036,64'hbf8d789c65167b66,
64'hcfc760b23833fa1a,64'hb6fc7a16c22e12db,64'h080b0692c120ee99,64'hb2a043752e8cf9ac,
64'hf22e934cec4d6a38,64'h2048fb04e1c0ae0f,64'h5a869e56d8353102,64'hc462328a529393c6,
64'h8214c5468193200c,64'h4bb1b026df98507d,64'hb4d653baa1f71121,64'ha6b394600e9ca35c,
64'h523bc9c3a8f0babb,64'hcbe38ac4345a71ee,64'h3f18c5f88f19f9fd,64'h52a870c4a011519b,
64'hbfe52ed67447f0e7,64'h3d7de67bea699f2b,64'h1c4e4d003ae61ab1,64'h0001000000000000,
64'ha7ea89586a5da9ce,64'h47c9bfee53a9b717,64'h2d3e749c32068452,64'h6564115e40c74369,
64'h01b38dbebdfa6116,64'h3a2d221e921a4d98,64'h566d77bf6373f366,64'h4bd6bb172e15d48c,
64'h7c37c1b35c27f705,64'h3642c4ee4d2e8c21,64'hcc11aab18ff446c8,64'h1e55b052fdb2e2c5,
64'he03c87747add3ecb,64'h05a66beefeca82ae,64'ha3895b400ec4b7d2,64'hc5c61f8349dd5fc6,
64'h3fe2eec3d33d2a6a,64'haeeb014cf9ddcd47,64'h777f917510a2cb72,64'h021f33dd513f8478,
64'h130718e613273091,64'hdc494cac0e52c375,64'h8eee94b90493fead,64'h8efb82c7d51bbde2,
64'hcb2fe38986336f49,64'h655c6bcd7533cc56,64'h484af27ff41fc8ce,64'hd317b839eae41235,
64'h5c2f2e47bb2809ef,64'hfb5dd0ce3b6df5c0,64'h7970df1e86ad2745,64'hffffffbeffc00041,
64'h4125e148fa9d3108,64'heec6e8cf5d74311c,64'h5a8943361a4d1411,64'hda274f509b042735,
64'h0ee85a03cf04b7b4,64'hfee0541488329da5,64'hed0e610eae3ad206,64'hbf96a7c861ef0ce4,
64'h9d07a93226f0dfda,64'h10022bde1b794cde,64'h507ab0504cb6a607,64'h57f1af134ca2cf6d,
64'hd9f8ec1587067f44,64'hb6df8f423845c25c,64'he10160d178241dd4,64'h9654086e25d19f36,
64'h1e45d2699d89ad47,64'h24091f607c3815c2,64'hcb50d3ca1b06a621,64'h588c46510a527279,
64'h904298a850326402,64'h697636047bf30a10,64'hf69aca76743ee225,64'h94d6728b81d3946c,
64'haa477937d51e1758,64'h597c7158468b4e3e,64'h67e318beb1e33f40,64'haa550e17f4022a34,
64'h37fca5daae88fe1d,64'ha7afbccedd4d33e6,64'he389c99f275cc357,64'h0000200000000000,
64'h54fd512acd4bb53a,64'h28f937fdaa7536e3,64'hc5a7ce92c640d08b,64'hecac822ae818e86e,
64'h403671b797bf4c23,64'h0745a443d24349b3,64'h4acdaef7ac6e7e6d,64'h897ad76265c2ba92,
64'h6f86f8360b84fee1,64'he6c8589ce9a5d185,64'h1982355631fe88d9,64'h63cab609ffb65c59,
64'hbc0790edef5ba7da,64'h40b4cd7d9fd95056,64'hd4712b6741d896fb,64'h58b8c3f0293babf9,
64'hc7fc5dd7ba67a54e,64'h35dd60297f3bb9a9,64'hceeff22de214596f,64'h0043e67baa27f08f,
64'he260e31be264e613,64'h7b89299521ca586f,64'h71ddd296c0927fd6,64'hd1df70583aa377bd,
64'hf965fc7050c66dea,64'h4cab8d796ea6798b,64'h49095e4fbe83f91a,64'h7a62f706dd5c8247,
64'h2b85e5c8d765013e,64'h1f6bba19c76dbeb8,64'h6f2e1be370d5a4e9,64'hfffffff6fff80009,
64'h0824bc291f53a621,64'h9dd8dd196bae8624,64'heb512865e349a283,64'h7b44e9e9b36084e7,
64'h81dd0b3ff9e096f7,64'h7fdc0a82310653b5,64'h5da1cc2195c75a41,64'h97f2d4f88c3de19d,
64'hd3a0f52584de1bfc,64'h4200457b836f299c,64'h2a0f5609e996d4c1,64'h6afe35e2099459ee,
64'h9b3f1d8230e0cfe9,64'h96dbf1e7c708b84c,64'h9c202c19af0483bb,64'h52ca810d84ba33e7,
64'h23c8ba4d13b135a9,64'hc48123eb4f8702b9,64'hf96a1a786360d4c5,64'heb1188c9414a4e50,
64'hd20853144a064c81,64'h0d2ec6c08f7e6142,64'h7ed3594e6e87dc45,64'h929ace50f03a728e,
64'h1548ef26faa3c2eb,64'h4b2f8e2ac8d169c8,64'h0cfc6317d63c67e8,64'h954aa1c27e804547,
64'h66ff94baf5d11fc4,64'h54f5f7999ba9a67d,64'h3c713933c4eb986b,64'h0000040000000000,
64'hca9faa2499a976a8,64'ha51f26ff154ea6dd,64'hb8b4f9d1b8c81a12,64'h5d9590451d031d0e,
64'ha806ce3652f7e985,64'ha0e8b487da486937,64'h6959b5de958dcfce,64'hd12f5aeb8cb85753,
64'hedf0df05e1709fdd,64'h7cd90b133d34ba31,64'he33046a9e63fd11c,64'hec7956c05ff6cb8c,
64'hd780f21cfdeb74fc,64'h481699af73fb2a0b,64'hba8e256c483b12e0,64'heb17187d25277580,
64'h58ff8bbab74cf4aa,64'he6bbac044fe77736,64'h39ddfe459c428b2e,64'h20087ccf5544fe12,
64'hbc4c1c62dc4c9cc3,64'h2f71253284394b0e,64'h4e3bba5298124ffb,64'h7a3bee0aa7546ef8,
64'hdf2cbf8d4a18cdbe,64'ha99571ae8dd4cf32,64'hc9212bc937d07f24,64'h2f4c5ee0bbab9049,
64'h4570bcb8daeca028,64'h03ed774338edb7d7,64'hede5c37b8e1ab49e,64'hfffffffdffff0002,
64'he104978443ea74c5,64'h93bb1ba2ad75d0c5,64'hbd6a250c1c693451,64'h2f689d3d166c109d,
64'h303ba167df3c12df,64'h6ffb814fe620ca77,64'hebb4398352b8eb49,64'h72fe5a9eb187bc34,
64'h9a741ea4309bc380,64'h884008aef06de534,64'he541eac05d32da99,64'h4d5fc6bc01328b3e,
64'hf367e3af661c19fe,64'h92db7e3c78e1170a,64'hb384058295e09078,64'h2a5950219097467d,
64'he4791748c27626b6,64'hf890247c89f0e058,64'h7f2d434eac6c1a99,64'h1d623119282949ca,
64'hfa410a61a940c991,64'hc1a5d8d751efcc29,64'h6fda6b296dd0fb89,64'h525359c9de074e52,
64'ha2a91de43f54785e,64'h0965f1c5591a2d39,64'h019f8c62fac78cfd,64'h32a954382fd008a9,
64'h8cdff296deba23f9,64'h6a9ebef2d37534d0,64'ha78e2725d89d730e,64'h0000008000000000,
64'h1953f54493352ed5,64'h74a3e4df82a9d4dc,64'hd7169f3977190343,64'h4bb2b20863a063a2,
64'h7500d9c66a5efd31,64'h341d1690db490d27,64'h4d2b36bb92b1b9fa,64'hba25eb5cd1970aeb,
64'h7dbe1be05c2e13fc,64'hef9b216187a69747,64'h9c6608d4bcc7fa24,64'h9d8f2ad78bfed972,
64'h9af01e431fbd6ea0,64'ha902d3354e7f6542,64'h1751c4ad8907625c,64'h1d62e30fa4a4eeb0,
64'hcb1ff17696e99e96,64'h5cd7758049fceee7,64'h473bbfc873885166,64'hc4010f992aa89fc3,
64'hb789838bbb899399,64'h45ee24a610872962,64'ha9c77749b3024a00,64'h0f477dc154ea8ddf,
64'h5be597f1694319b8,64'hd532ae3511ba99e7,64'h99242578a6fa0fe5,64'he5e98bdb3775720a,
64'h08ae17971b5d9405,64'h207daee8471db6fb,64'h5dbcb86f31c35694,64'hdffffffeffffe001,
64'h7c2092f0287d4e99,64'h72776373f5aeba19,64'hf7ad44a0a38d268b,64'h65ed13a742cd8214,
64'h2607742cdbe7825c,64'h2dff7029dcc4194f,64'hfd76872f8a571d6a,64'h8e5fcb535630f787,
64'h134e83d486137870,64'h910801155e0dbca7,64'hfca83d572ba65b54,64'h49abf8d740265168,
64'h5e6cfc75acc38340,64'hd25b6fc6cf1c22e2,64'h167080b052bc120f,64'h654b2a03d212e8d0,
64'h5c8f22e8d84ec4d7,64'h1f12048f913e1c0b,64'hefe5a868f58d8354,64'hc3ac46226505293a,
64'hff48214b55281933,64'hf834bb1a0a3df986,64'hedfb4d644dba1f72,64'hca4a6b387bc0e9cb,
64'h545523bc47ea8f0c,64'he12cbe37cb2345a8,64'h6033f18bff58f1a0,64'he6552a8625fa0116,
64'hf19bfe51fbd74480,64'h0d53d7de5a6ea69a,64'h54f1c4e47b13ae62,64'h0000001000000000,
64'h632a7ea83266a5db,64'h8e947c9b70553a9c,64'hbae2d3e68ee32069,64'hc97656404c740c75,
64'heea01b37ed4bdfa7,64'h2683a2d1fb6921a5,64'hc9a566d6b2563740,64'hb744bd6afa32e15e,
64'h8fb7c37b8b85c280,64'h3df3642c10f4d2e9,64'h938cc11a1798ff45,64'hd3b1e55a317fdb2f,
64'h135e03c863f7add4,64'hd5205a65e9cfeca9,64'h82ea38953120ec4c,64'h03ac5c61f4949dd6,
64'h5963fe2e92dd33d3,64'h2b9aeeafe93f9ddd,64'h48e777f8ce710a2d,64'hb88021f2855513f9,
64'hf6f1307097713274,64'hc8bdc4940210e52d,64'h1538eee936604940,64'h21e8efb80a9d51bc,
64'h0b7cb2fe2d286337,64'h3aa655c68237533d,64'h732484aeb4df41fd,64'hdcbd317aa6eeae42,
64'h6115c2f2836bb281,64'ha40fb5dc68e3b6e0,64'h8bb7970d66386ad3,64'hfbfffffefffffc01,
64'hef84125d250fa9d4,64'hee4eec6d9eb5d744,64'hbef5a8937471a4d2,64'h8cbda2746859b043,
64'h84c0ee851b7cf04c,64'h25bfee051b98832a,64'hdfaed0e5314ae3ae,64'h31cbf96a4ac61ef1,
64'h0269d07a90c26f0e,64'h322100228bc1b795,64'h9f9507aa6574cb6b,64'h09357f1ae804ca2d,
64'h0bcd9f8eb5987068,64'hda4b6df819e3845d,64'h22ce1015ea578242,64'h0ca965407a425d1a,
64'h2b91e45cfb09d89b,64'ha3e240915227c382,64'h9dfcb50c9eb1b06b,64'hd87588c38ca0a528,
64'hbfe90428caa50327,64'h5f0697630147bf31,64'hddbf69abc9b743ef,64'hb9494d666f781d3a,
64'h8a8aa47708fd51e2,64'h1c2597c6f96468b5,64'h0c067e317feb1e34,64'h5ccaa55084bf4023,
64'h1e337fca3f7ae890,64'hc1aa7afb0b4dd4d4,64'hca9e389bcf6275cd,64'h0000000200000000,
64'hac654fd4664cd4bc,64'h91d28f92ee0aa754,64'hf75c5a7bf1dc640e,64'h792ecac7a98e818f,
64'h3dd40366dda97bf5,64'h64d07459df6d2435,64'h1934acdad64ac6e8,64'h56e897ad1f465c2c,
64'h11f6f86f7170b850,64'he7be6c84a21e9a5e,64'h72719822e2f31fe9,64'h3a763cab262ffb66,
64'h826bc0788c7ef5bb,64'hfaa40b4bdd39fd96,64'h905d471226241d8a,64'h40758b8bfe9293bb,
64'hab2c7fc5325ba67b,64'h65735dd59d27f3bc,64'h691ceefeb9ce2146,64'hf710043d70aaa280,
64'h9ede260d92ee264f,64'h7917b89220421ca6,64'h02a71ddd26cc0928,64'h843d1df68153aa38,
64'h216f965fa5a50c67,64'h6754cab87046ea68,64'h6e649095769be840,64'hdb97a62e94ddd5c9,
64'hec22b85d706d7651,64'h1481f6bb8d1c76dc,64'hb176f2e10cc70d5b,64'hff7ffffeffffff81,
64'h9df0824b24a1f53b,64'h9dc9dd8d33d6bae9,64'hd7deb511ae8e349b,64'hb197b44ded0b3609,
64'h90981dd0236f9e0a,64'hc4b7fdbfe3731066,64'h5bf5da1c66295c76,64'he6397f2c6958c3df,
64'h404d3a0f12184de2,64'h66442003f17836f3,64'hb3f2a0f4acae996e,64'h6126afe2fd009946,
64'h0179b3f1d6b30e0d,64'h7b496dbea33c708c,64'hc459c201fd4af049,64'hc1952ca74f484ba4,
64'ha5723c8aff613b14,64'hd47c48116a44f871,64'hb3bf96a0f3d6360e,64'h1b0eb118719414a5,
64'h37fd2084f954a065,64'hebe0d2eb8028f7e7,64'h3bb7ed355936e87e,64'hd72929ac0def03a8,
64'hd151548e211faa3d,64'h6384b2f87f2c8d17,64'h8180cfc5affd63c7,64'hab9954a97097e805,
64'h03c66ff947ef5d12,64'h98354f5ee169ba9b,64'h7953c71319ec4eba,64'h0000000040000000,
64'h958ca9fa0cc99a98,64'h923a51f1ddc154eb,64'h5eeb8b4f3e3b8c82,64'h2f25d958d531d032,
64'h67ba806c7bb52f7f,64'h6c9a0e8adbeda487,64'h0326959b5ac958dd,64'h8add12f523e8cb86,
64'h023edf0dee2e170a,64'h5cf7cd905443d34c,64'hee4e33037c5e63fe,64'h474ec79524c5ff6d,
64'hb04d780e718fdeb8,64'h5f5481693ba73fb3,64'hd20ba8e184c483b2,64'ha80eb170dfd25278,
64'hb5658ff8064b74d0,64'h8cae6bba33a4fe78,64'h4d239ddf9739c429,64'h1ee20087ae155450,
64'h33dbc4c1925dc4ca,64'h4f22f71204084395,64'h0054e3bba4d98125,64'h1087a3bed02a7547,
64'h242df2cbd4b4a18d,64'h0cea99570e08dd4d,64'h0dcc9212aed37d08,64'hfb72f4c4f29bbaba,
64'hfd84570ace0daecb,64'h82903ed6f1a38edc,64'hb62ede5b8198e1ac,64'hffeffffefffffff1,
64'hb3be1048c4943ea8,64'hf3b93bb0c67ad75e,64'hbafbd6a195d1c694,64'hf632f688dda166c2,
64'hd21303b9446df3c2,64'h5896ffb7bc6e620d,64'h4b7ebb434cc52b8f,64'h3cc72fe56d2b187c,
64'hc809a741224309bd,64'hacc883ffde2f06df,64'h567e541e5595d32e,64'h4c24d5fc1fa01329,
64'h602f367ddad661c2,64'h8f692db754678e12,64'hf88b383f5fa95e0a,64'h9832a59469e90975,
64'h94ae4790dfec2763,64'hfa8f89014d489f0f,64'h5677f2d3de7ac6c2,64'h6361d622ae328295,
64'h66ffa4103f2a940d,64'h3d7c1a5d50051efd,64'h4776fda66b26dd10,64'h1ae5253581bde075,
64'h7a2a2a916423f548,64'h2c70965eefe591a3,64'h303019f895ffac79,64'h75732a94ce12fd01,
64'hc078cdfe68fdeba3,64'hb306a9eb3c2d3754,64'hcf2a78e1a33d89d8,64'h0000000008000000,
64'h12b1953f41993353,64'hb2474a3d9bb82a9e,64'hcbdd716927c77191,64'hc5e4bb2a5aa63a07,
64'h2cf7500d6f76a5f0,64'h2d9341d13b7db491,64'h6064d2b30b592b1c,64'h515ba25e647d1971,
64'hc047dbe0fdc5c2e2,64'h8b9ef9b18a887a6a,64'h5dc9c6602f8bcc80,64'h68e9d8f24498bfee,
64'h1609af01ce31fbd7,64'habea902c8774e7f7,64'hda41751b70989077,64'h1501d62e1bfa4a4f,
64'h16acb1ff00c96e9a,64'h1195cd7746749fcf,64'he9a473bb12e73886,64'h03dc4010f5c2aa8a,
64'hc67b7897724bb89a,64'h69e45ee1e0810873,64'h600a9c77149b3025,64'h2210f477ba054ea9,
64'h6485be591a969432,64'h619d532a81c11baa,64'h01b9924255da6fa1,64'hdf6e5e97de537758,
64'hbfb08ae0b9c1b5da,64'h905207da5e3471dc,64'h96c5dbcaf0331c36,64'hfffdfffeffffffff,
64'h1677c209189287d5,64'h5e772775d8cf5aec,64'h975f7ad3b2ba38d3,64'hdec65ed05bb42cd9,
64'hda426076688dbe79,64'h6b12dff6978dcc42,64'h296fd7684998a572,64'h8798e5fc2da56310,
64'h790134e7c4486138,64'h3599107fdbc5e0dc,64'h4acfca838ab2ba66,64'he9849abea3f40266,
64'hcc05e6cefb5acc39,64'hd1ed25b62a8cf1c3,64'hdf1167072bf52bc2,64'h730654b22d3d212f,
64'hb295c8f17bfd84ed,64'h3f51f12009a913e2,64'hcacefe59bbcf58d9,64'h6c6c3ac3f5c65053,
64'h6cdff481a7e55282,64'h67af834b4a00a3e0,64'h08eedfb4cd64dba2,64'h635ca4a65037bc0f,
64'h0f4545522c847ea9,64'ha58e12cb3dfcb235,64'he606033e32bff590,64'heeae6551b9c25fa1,
64'hb80f19bf2d1fbd75,64'h9660d53ce785a6eb,64'h19e54f1c3467b13b,64'h0000000001000000,
64'ha25632a74833266b,64'h5648e94773770554,64'hf97bae2c44f8ee33,64'h38bc97652b54c741,
64'h059eea01adeed4be,64'he5b26839476fb693,64'h8c0c9a55e16b2564,64'hea2b744aec8fa32f,
64'hd808fb7b5fb8b85d,64'hd173df3571510f4e,64'h0bb938cc05f17990,64'h4d1d3b1e089317fe,
64'h22c135e019c63f7b,64'h357d520570ee9cff,64'h3b482ea34e13120f,64'h22a03ac5a37f494a,
64'hc2d5963f20192dd4,64'h2232b9aec8ce93fa,64'h5d348e77225ce711,64'hc07b88015eb85552,
64'hd8cf6f122e497714,64'had3c8bdb9c10210f,64'h6c01538e82936605,64'he4421e8e1740a9d6,
64'hcc90b7ca6352d287,64'hcc33aa6490382376,64'he03732476abb4df5,64'h1bedcbd2fbca6eeb,
64'hd7f6115b573836bc,64'h920a40facbc68e3c,64'h52d8bb791e066387,64'h3fffbfffc0000000,
64'h62cef840c31250fb,64'h8bcee4ee3b19eb5e,64'hb2ebef59d657471b,64'hfbd8cbd92b76859c,
64'hfb484c0ded11b7d0,64'hcd625bfe12f1b989,64'hc52dfaec493314af,64'h10f31cbf85b4ac62,
64'h0f20269cf8890c27,64'h86b3220f7b78bc1c,64'h4959f9503156574d,64'h5d309357947e804d,
64'hf980bcd8ff6b5988,64'hba3da4b625519e39,64'hdbe22ce0257ea579,64'h2e60ca9625a7a426,
64'h7652b91dcf7fb09e,64'hc7ea3e234135227d,64'hf959dfca5779eb1c,64'had8d8757deb8ca0b,
64'hcd9bfe8f74fcaa51,64'h0cf5f0696940147c,64'hc11ddbf5d9ac9b75,64'h2c6b9494aa06f782,
64'he1e8a8a965908fd6,64'h74b1c25907bf9647,64'h1cc0c067c657feb2,64'hfdd5cca957384bf5,
64'h7701e33785a3f7af,64'hb2cc1aa6fcf0b4de,64'ha33ca9e2e68cf628,64'h0000000000200000,
64'hb44ac654490664ce,64'h8ac91d286e6ee0ab,64'hbf2f75c4e89f1dc7,64'he71792ebc56a98e9,
64'h40b3dd3ff5bdda98,64'hbcb64d0688edf6d3,64'h9181934a3c2d64ad,64'h3d456e893d91f466,
64'h7b011f6f0bf7170c,64'h5a2e7be66e2a21ea,64'h0177271980be2f32,64'h49a3a76381126300,
64'ha45826bb6338c7f0,64'h26afaa408e1dd3a0,64'h276905d449c26242,64'hc4540757f46fe92a,
64'h985ab2c7640325bb,64'hc44657351919d280,64'heba691ce044b9ce3,64'hd80f70ff6bd70aab,
64'h9b19ede1c5c92ee3,64'h35a7917b53820422,64'h6d802a7170526cc1,64'h5c8843d182e8153b,
64'h399216f92c6a5a51,64'h5986754c5207046f,64'h7c06e6488d5769bf,64'ha37db979bf794dde,
64'h9afec22aeae706d8,64'h9241481ed978d1c8,64'h2a5b176f03c0cc71,64'h07fff7fff8000000,
64'hac59df0778624a20,64'h5179dc9d87633d6c,64'hb65d7dea9acae8e4,64'h9f7b197aa56ed0b4,
64'h1f690981bda236fa,64'hf9ac4b7ee25e3732,64'h38a5bf5d69266296,64'hc21e639730b6958d,
64'h21e404d37f112185,64'h90d664416f6f1784,64'h692b3f29a62acaea,64'h6ba6126a928fd00a,
64'h1f30179b1fed6b31,64'hf747b495e4aa33c8,64'hfb7c459b24afd4b0,64'h45cc195284b4f485,
64'h4eca572379eff614,64'h78fd47c40826a450,64'h9f2b3bf8caef3d64,64'hb5b1b0ea5bd71942,
64'hf9b37fd10e9f954b,64'h819ebe0cad280290,64'h7823bb7e5b35936f,64'hc58d7291d540def1,
64'h5c3d1514ecb211fb,64'h2e96384b00f7f2c9,64'hc398180c38caffd7,64'h7fbab994cae7097f,
64'h2ee03c66d0b47ef6,64'h565983549f9e169c,64'h1467953c5cd19ec5,64'h0000000000040000,
64'h568958ca4920cc9a,64'hb15923a46dcddc16,64'h37e5eeb87d13e3b9,64'hfce2f25c98ad531e,
64'h08167ba7feb7bb53,64'hb796c9a0311dbedb,64'h72303268e785ac96,64'h47a8add0e7b23e8d,
64'h8f6023ed617ee2e2,64'hcb45cf7c0dc5443e,64'hc02ee4e27017c5e7,64'h093474ec70224c60,
64'h148b04d76c6718fe,64'h04d5f54811c3ba74,64'hc4ed20b9c9384c49,64'hd88a80ea3e8dfd26,
64'hb30b56584c8064b8,64'h1888cae6a3233a50,64'hbd74d2392089739d,64'hbb01ee1f4d7ae156,
64'hb3633dbb98b925dd,64'hc6b4f22eaa704085,64'hedb0054d4e0a4d99,64'hab910879905d02a8,
64'he73242de458d4b4b,64'h2b30cea96a40e08e,64'h2f80dcc8f1aaed38,64'h546fb72ef7ef29bc,
64'h135fd8455d5ce0db,64'h12482903db2f1a39,64'he54b62ed0078198f,64'h00fffeffff000000,
64'h158b3be0ef0c4944,64'h8a2f3b9330ec67ae,64'h96cbafbcd3595d1d,64'h93ef632ed4adda17,
64'hc3ed212f77b446e0,64'hdf35896f1c4bc6e7,64'h4714b7eb6d24cc53,64'h7843cc728616d2b2,
64'h643c809a0fe22431,64'h921acc87adede2f1,64'hcd2567e474c5595e,64'hcd74c24c9251fa02,
64'he3e602f283fdad67,64'h1ee8f692bc954679,64'h1f6f88b36495fa96,64'h68b98329f0969e91,
64'h89d94ae3ef3dfec3,64'h0f1fa8f88104d48a,64'h93e5677e995de7ad,64'hd6b6361c8b7ae329,
64'hbf366ff981d3f2aa,64'h1033d7c195a50052,64'h2f04776fab66b26e,64'hf8b1ae515aa81bdf,
64'hab87a2a1fd964240,64'he5d2c708801efe5a,64'h3873030167195ffb,64'h2ff75732795ce130,
64'h45dc078c9a168fdf,64'h8acb306a13f3c2d4,64'h628cf2a72b9a33d9,64'h0000000000008000,
64'hcad12b1889241994,64'h562b24744db9bb83,64'he6fcbdd62fa27c78,64'h5f9c5e4b5315aa64,
64'ha102cf745fd6f76b,64'hb6f2d9336623b7dc,64'h4e46064cdcf0b593,64'h68f515b9bcf647d2,
64'hd1ec047cec2fdc5d,64'h5968b9ef41b8a888,64'h3805dc9c2e02f8bd,64'h01268e9d8e04498c,
64'h4291609aad8ce320,64'h809abea88238774f,64'hf89da4165927098a,64'h5b11501d07d1bfa5,
64'h16616acb09900c97,64'h0311195cd464674a,64'h77ae9a46c4112e74,64'h57603dc3a9af5c2b,
64'h766c67b7131724bc,64'h78d69e45754e0811,64'hfdb600a8c9c149b4,64'h1572210f320ba055,
64'hbce6485b28b1a96a,64'h456619d4ed481c12,64'h05f01b991e355da7,64'h8a8df6e55efde538,
64'ha26bfb080bab9c1c,64'he249051f9b65e348,64'h3ca96c5d800f0332,64'h001fffdfffe00000,
64'h82b1677b9de18929,64'h5145e772261d8cf6,64'h72d975f73a6b2ba4,64'h327dec65ba95bb43,
64'h187da425eef688dc,64'h3be6b12dc38978dd,64'ha8e296fccda4998b,64'hcf08798d90c2da57,
64'hec87901261fc4487,64'hf243599015bdbc5f,64'h59a4acfc4e98ab2c,64'hd9ae9848d24a3f41,
64'h3c7cc05e307fb5ad,64'he3dd1ed17792a8d0,64'h43edf1162c92bf53,64'hed1730645e12d3d3,
64'hb13b295bdde7bfd9,64'hc1e3f51e50209a92,64'h727cacef732bbcf6,64'hfad6c6c2b16f5c66,
64'hd7e6cdfe703a7e56,64'hc2067af772b4a00b,64'h45e08eedb56cd64e,64'h3f1635ca0b55037c,
64'h1570f4543fb2c848,64'hdcba58e05003dfcc,64'ha70e605f8ce32c00,64'h05feeae64f2b9c26,
64'h28bb80f17342d1fc,64'h9159660cc27e785b,64'hec519e540573467c,64'h0000000000001000,
64'h995a256291248333,64'haac5648de9b73771,64'h1cdf97bac5f44f8f,64'h8bf38bc8ea62b54d,
64'hb42059edebfadeee,64'h96de5b25ecc476fc,64'ha9c8c0c8fb9e16b3,64'hcd1ea2b6779ec8fb,
64'h7a3d808f3d85fb8c,64'h0b2d173de8371511,64'h6700bb9325c05f18,64'h8024d1d331c08932,
64'h08522c1355b19c64,64'h301357d4f0470eea,64'hdf13b4820b24e132,64'h6b622a0340fa37f5,
64'h22cc2d5941320193,64'hc062232ada8c8cea,64'h8ef5d348588225cf,64'haaec07b7d535eb86,
64'h8ecd8cf66262e498,64'hef1ad3c7cea9c103,64'h9fb6c01499382937,64'h62ae44218641740b,
64'hd79cc90aa516352e,64'hc8acc339dda90383,64'h20be037303c6abb5,64'h1151bedcabdfbca7,
64'h944d7f6081757384,64'h1c4920a3f36cbc69,64'hc7952d8af001e067,64'h0003fffbfffc0000,
64'hf0562cee93bc3126,64'h4a28bcee04c3b19f,64'h8e5b2ebe674d6575,64'ha64fbd8c1752b769,
64'h830fb4843dded11c,64'h677cd62558712f1c,64'hb51c52def9b49332,64'h39e10f3192185b4b,
64'h3d90f2022c3f8891,64'h3e486b31e2b7b78c,64'h8b34959f09d31566,64'hfb35d3083a4947e9,
64'h678f980b660ff6b6,64'h1c7ba3da2ef2551a,64'ha87dbe22259257eb,64'hbda2e60bebc25a7b,
64'hf627652a9bbcf7fc,64'hd83c7ea30a041353,64'h4e4f959dae65779f,64'h5f5ad8d8162deb8d,
64'h5afcd9bf8e074fcb,64'hb840cf5e4e569402,64'h48bc11dd76ad9aca,64'h87e2c6b8c16aa070,
64'h02ae1e8a87f65909,64'h9b974b1b8a007bfa,64'h14e1cc0bf19c6580,64'h40bfdd5c89e57385,
64'h8517701dae685a40,64'hb22b2cc0f84fcf0c,64'h9d8a33ca00ae68d0,64'h0000000000000200,
64'hb32b44abb2249067,64'hf558ac90dd36e6ef,64'h239bf2f738be89f2,64'h717e7178bd4c56aa,
64'h56840b3d7d7f5bde,64'h92dbcb643d988ee0,64'hb53918187f73c2d7,64'hb9a3d4562ef3d920,
64'h8f47b01167b0bf72,64'he165a2e6dd06e2a3,64'h0ce0177264b80be3,64'hd0049a39a6381127,
64'h810a4581eab6338d,64'hc6026af9de08e1de,64'hdbe2768f81649c27,64'h6d6c4540081f46ff,
64'ha45985aa88264033,64'hd80c44649b51919e,64'h31deba68eb1044ba,64'h555d80f6baa6bd71,
64'h11d9b19ecc4c5c93,64'hbde35a7859d53821,64'h33f6d80273270527,64'hac55c88390c82e82,
64'h5af3992114a2c6a6,64'hb91598669bb52071,64'h6417c06e0078d577,64'h222a37db757bf795,
64'h9289afeb902eae71,64'he38924139e6d978e,64'h38f2a5b13e003c0d,64'h00007fff7fff8000,
64'h5e0ac59d92778625,64'h2945179da0987634,64'h71cb65d76ce9acaf,64'hf4c9f7b0a2ea56ee,
64'h9061f69007bbda24,64'h8cef9ac42b0e25e4,64'hd6a38a5b1f369267,64'ha73c21e592430b6a,
64'he7b21e3f6587f113,64'h87c90d65bc56f6f2,64'h516692b3a13a62ad,64'hff66ba60274928fe,
64'h4cf1f3012cc1fed7,64'hc38f747a85de4aa4,64'hb50fb7c3a4b24afe,64'hb7b45cc0dd784b50,
64'h9ec4eca4d3779f00,64'hbb078fd3c140826b,64'h29c9f2b395ccaef4,64'h6beb5b1aa2c5bd72,
64'hab5f9b3751c0e9fa,64'hd70819eb09cad281,64'hc917823aeed5b35a,64'h10fc58d7182d540e,
64'he055c3d070fecb22,64'hd372e962b1400f80,64'h029c39817e338cb0,64'h6817fbab313cae71,
64'h10a2ee03b5cd0b48,64'h964565979f09f9e2,64'h13b146794015cd1a,64'h0000000000000040,
64'h366568955644920d,64'h3eab1591fba6dcde,64'hc4737e5e2717d13f,64'hce2fce2e57a98ad6,
64'h4ad081676fafeb7c,64'h125b796c87b311dc,64'h36a72302efee785b,64'h17347a8ac5de7b24,
64'hd1e8f6016cf617ef,64'hbc2cb45c3ba0dc55,64'ha19c02edac97017d,64'h3a00934714c70225,
64'h702148afdd56c672,64'h58c04d5efbc11c3c,64'h3b7c4ed1d02c9385,64'h2dad88a7e103e8e0,
64'hb48b30b4b104c807,64'h5b01888c536a3234,64'hc63bd74c5d620898,64'heaabb01df754d7af,
64'ha23b363339898b93,64'hf7bc6b4e2b3aa705,64'h267edb002e64e0a5,64'hd58ab90fb21905d1,
64'h4b5e7323e29458d5,64'hf722b30bf376a40f,64'h2c82f80da00f1aaf,64'h644546fb0eaf7ef3,
64'hf25135fc9205d5cf,64'h5c71248233cdb2f2,64'h671e54b5c7c00782,64'h00000fffeffff000,
64'h6bc158b3524ef0c5,64'h8528a2f334130ec7,64'h2e396cbacd9d3596,64'h5e993ef5d45d4ade,
64'h920c3ed180f77b45,64'h919df3580561c4bd,64'h3ad4714b43e6d24d,64'hd4e7843bf248616e,
64'hbcf643c74cb0fe23,64'hd0f921abf78adedf,64'h6a2cd25614274c56,64'h5fecd74bc4e92520,
64'h299e3e6005983fdb,64'h9871ee8ed0bbc955,64'h56a1f6f834964960,64'h16f68b981baf096a,
64'h13d89d949a6ef3e0,64'hb760f1f9d828104e,64'h85393e55f2b995df,64'hcd7d6b629458b7af,
64'hd56bf3662a381d40,64'hfae1033c81395a51,64'hd922f0469ddab66c,64'h421f8b1aa305aa82,
64'hdc0ab8794e1fd965,64'h1a6e5d2c562801f0,64'h005387302fc67196,64'hed02ff74862795cf,
64'h02145dc076b9a169,64'hd2c8acb233e13f3d,64'hc27628ce6802b9a4,64'h0000000000000008,
64'h66ccad124ac89242,64'h47d562b1ff74db9c,64'h388e6fcba4e2fa28,64'h59c5f9c58af5315b,
64'h895a102c6df5fd70,64'h824b6f2d10f6623c,64'ha6d4e45fbdfdcf0c,64'h82e68f50d8bbcf65,
64'h3a3d1ec00d9ec2fe,64'h7785968b27741b8b,64'h7433805d5592e030,64'h674012688298e045,
64'hce0429153baad8cf,64'h8b1809ab5f782388,64'h676f89d9da059271,64'h05b5b114fc207d1c,
64'h3691661676209901,64'h8b6031110a6d4647,64'h18c77ae98bac4113,64'h3d5576039eea9af6,
64'hb44766c5c7313173,64'h7ef78d69656754e1,64'h64cfdb5fa5cc9c15,64'hfab15721164320bb,
64'h696bce641c528b1b,64'h3ee456615e6ed482,64'h25905f019401e356,64'hac88a8dec1d5efdf,
64'h3e4a26bf7240baba,64'hcb8e248f8679b65f,64'hcce3ca95f8f800f1,64'h000001fffdfffe00,
64'h6d782b160a49de19,64'h30a5145e468261d9,64'h45c72d9719b3a6b3,64'h4bd327de7a8ba95c,
64'h724187d9d01eef69,64'h7233be6aa0ac3898,64'h675a8e29087cda4a,64'h5a9cf0873e490c2e,
64'hb79ec87849961fc5,64'h3a1f24355ef15bdc,64'h4d459a4a8284e98b,64'h0bfd9ae9789d24a4,
64'ha533c7cb60b307fc,64'h730e3dd17a17792b,64'h0ad43edf0692c92c,64'hc2ded1724375e12e,
64'h027b13b2934dde7c,64'h56ec1e3efb05020a,64'h30a727ca9e5732bc,64'h39afad6c328b16f6,
64'h1aad7e6cc54703a8,64'hff5c2066b0272b4b,64'h9b245e0853bb56ce,64'hc843f1629460b551,
64'h7b81570ec9c3fb2d,64'h034dcba58ac5003e,64'h400a70e5c5f8ce33,64'h3da05fee70c4f2ba,
64'he0428bb72ed7342e,64'h7a591595e67c27e8,64'h984ec5194d005735,64'h0000000000000001
};
  //------------------------
  // 1024
  //------------------------
  localparam [2*1024-1:0][63:0] NTT_GF64_FWD_N1024_PHI_L = {
64'h88faac55bfee9b74,64'hab38bf38115ea62c,64'h90496de5221ecc48,64'h705cd1e9bb1779ed,
64'haef0b2d0c4ee8372,64'h6ce8024cb0531c09,64'h116301356bef0471,64'h80b6b6221f840fa4,
64'h316c0622014da8c9,64'h47aaaec033dd535f,64'hefdef1ac4cacea9d,64'hbf562ae382c86418,
64'hc7dc8acb6bcdda91,64'h3591151bb83abdfc,64'h3971c491d0cf36cc,64'h0000003fffbfffc0,
64'he614a28ae8d04c3c,64'h897a64fb4f51752c,64'h0e4677cd54158713,64'h4b539e10a7c92186,
64'h8743e4862bde2b7c,64'h817fb35caf13a495,64'hae61c7b98f42ef26,64'h585bda2e086ebc26,
64'hcadd83c71f60a042,64'h4735f5ad465162df,64'hbfeb840c3604e56a,64'hf9087e2b728c16ab,
64'h4069b9747158a008,64'hc7b40bfd0e189e58,64'h0f4b22b2bccf84fd,64'hdfffffff20000001,
64'h911f558a37fdd36f,64'h956717e6822bd4c6,64'h12092dbca443d989,64'h6e0b9a3cd762ef3e,
64'hd5de1659589dd06f,64'hed9d0048b60a6382,64'he22c6025cd7de08f,64'h9016d6c3c3f081f5,
64'he62d80c36029b51a,64'h28f555d7e67baa6c,64'h7dfbde3529959d54,64'h17eac55c70590c83,
64'hf8fb91588d79bb53,64'h86b222a2f70757c0,64'h872e3891ba19e6da,64'h00000007fff7fff8,
64'h9cc29450dd1a0988,64'h912f4c9ee9ea2ea6,64'ha1c8cef90a82b0e3,64'h496a73c1d4f92431,
64'h90e87c90457bc570,64'h702ff66b35e27493,64'h55cc38f6f1e85de5,64'h4b0b7b45810dd785,
64'hd95bb07823ec1409,64'h28e6beb588ca2c5c,64'hd7fd7080c6c09cae,64'hbf210fc4ce5182d6,
64'h080d372e8e2b1401,64'h18f6817fa1c313cb,64'h61e96455f799f0a0,64'hfbffffff04000001,
64'h3223eab126ffba6e,64'h52ace2fc90457a99,64'he24125b6b4887b32,64'h4dc173475aec5de8,
64'h3abbc2cb0b13ba0e,64'hddb3a00856c14c71,64'h3c458c0499afbc12,64'h7202dad8187e103f,
64'hdcc5b017ac0536a4,64'h851eaaba7ccf754e,64'h8fbf7bc62532b3ab,64'ha2fd58aaee0b2191,
64'hbf1f722a71af376b,64'h10d644545ee0eaf8,64'hd0e5c71177433cdc,64'h00000000fffeffff,
64'h1398528a1ba34131,64'h5225e9939d3d45d5,64'hb43919de8150561d,64'he92d4e775a9f2487,
64'h121d0f9208af78ae,64'hae05feccc6bc4e93,64'h6ab9871e7e3d0bbd,64'h69616f685021baf1,
64'hfb2b760e247d8282,64'h851cd7d63119458c,64'h5affae0fd8d81396,64'h57e421f859ca305b,
64'he101a6e4f1c56281,64'ha31ed02f5438627a,64'h0c3d2c8abef33e14,64'hff7fffff00800001,
64'h46447d55e4dff74e,64'hea559c5eb208af54,64'hdc4824b616910f67,64'h09b82e68eb5d8bbd,
64'h4757785921627742,64'hfbb674002ad8298f,64'hc788b17fd335f783,64'h2e405b5ae30fc208,
64'h9b98b6027580a6d5,64'h50a3d5570f99eeaa,64'hb1f7ef7824a65676,64'hf45fab147dc16433,
64'hb7e3ee44ae35e6ee,64'h021ac88a8bdc1d5f,64'h9a1cb8e1aee8679c,64'h1fffffffffffe000,
64'he2730a5063746827,64'h6a44bd3213a7a8bb,64'h7687233b702a0ac4,64'h3d25a9cecb53e491,
64'h4243a1f20115ef16,64'hb5c0bfd8f8d789d3,64'h6d5730e36fc7a178,64'hed2c2dec2a04375f,
64'hdf656ec1048fb051,64'h90a39afa462328b2,64'h4b5ff5c1bb1b0273,64'haafc843e6b39460c,
64'hfc2034dbbe38ac51,64'hd463da052a870c50,64'h8187a590d7de67c3,64'hffefffff00100001,
64'h48c88faa7c9bfeea,64'h9d4ab38b564115eb,64'h3b890496a2d221ed,64'h613705ccbd6bb178,
64'hc8eaef0a642c4ee9,64'h3f76ce7fe55b0532,64'hb8f1162f5a66bef1,64'h05c80b6b5c61f841,
64'h737316bfeeb014db,64'hca147aaa21f33dd6,64'h563efdeec494cacf,64'hbe8bf561efb82c87,
64'h56fc7dc855c6bcde,64'h20435911317b83ac,64'h9343971bb5dd0cf4,64'h03fffffffffffc00,
64'h3c4e6149ec6e8d05,64'had4897a5a274f518,64'h8ed0e466ee054159,64'he7a4b538f96a7c93,
64'h4848743e0022bde3,64'hb6b817fa7f1af13b,64'h0daae61c6df8f42f,64'h3da585bd654086ec,
64'hfbecadd74091f60b,64'hd214735e88c46517,64'ha96bfeb79763604f,64'h955f90874d6728c2,
64'hff84069a97c7158b,64'h1a8c7b40a550e18a,64'hb030f4b17afbccf9,64'hfffdffff00020001,
64'hc91911f48f937fde,64'hb3a95670cac822be,64'h67712092745a443e,64'h0c26e0b997ad762f,
64'hf91d5de06c8589de,64'hc7eed9cf3cab60a7,64'hf71e22c50b4cd7df,64'he0b9016c8b8c3f09,
64'hae6e62d75dd6029c,64'h59428f55043e67bb,64'h2ac7dfbdb892995a,64'h37d17eac1df70591,
64'h4adf8fb8cab8d79c,64'h84086b21a62f7076,64'h926872e2f6bba19f,64'h007fffffffffff80,
64'h6789cc28dd8dd1a1,64'h15a912f4b44e9ea3,64'hf1da1c8bfdc0a82c,64'hbcf496a67f2d4f93,
64'ha9090e87200457bd,64'hb6d702feafe35e28,64'h21b55cc36dbf1e86,64'h87b4b0b72ca810de,
64'hbf7d95ba48123ec2,64'h3a428e6bb1188ca3,64'h352d7fd6d2ec6c0a,64'hd2abf21029ace519,
64'hbff080d2b2f8e2b2,64'hc3518f6754aa1c32,64'hf6061e954f5f79a0,64'hffffbfff00004001,
64'h5923223e51f26ffc,64'h56752acdd9590458,64'h4cee24120e8b4888,64'h2184dc1712f5aec6,
64'h5f23abbbcd90b13c,64'h38fddb39c7956c15,64'h3ee3c45881699afc,64'hfc17202cb17187e2,
64'h95cdcc5a6bbac054,64'hab2851ea0087ccf8,64'hc558fbf6f712532c,64'he6fa2fd4a3bee0b3,
64'h895bf1f699571af4,64'h50810d63f4c5ee0f,64'h324d0e5c3ed77434,64'h000ffffffffffff0,
64'hecf139843bb1ba35,64'ha2b5225df689d3d5,64'h9e3b4390ffb81506,64'hb79e92d42fe5a9f3,
64'h752121d084008af8,64'h16dae05fd5fc6bc5,64'h4436ab982db7e3d1,64'h50f69616a595021c,
64'hd7efb2b6890247d9,64'ha74851ccd6231195,64'hc6a5affa1a5d8d82,64'hfa557e4125359ca4,
64'hd7fe1019965f1c57,64'hd86a31ec2a954387,64'h1ec0c3d2a9ebef34,64'hfffff7ff00000801,
64'h8b2464474a3e4e00,64'h0acea559bb2b208b,64'h099dc48241d16911,64'h44309b82a25eb5d9,
64'h8be47576f9b21628,64'h671fbb66d8f2ad83,64'h87dc788a902d3360,64'hdf82e404d62e30fd,
64'h92b9b98acd77580b,64'h15650a3d4010f99f,64'h98ab1f7e5ee24a66,64'hbcdf45f9f477dc17,
64'h912b7e3e532ae35f,64'h2a1021ac5e98bdc2,64'h8649a1cb07daee87,64'h0001fffffffffffe,
64'h7d9e273027763747,64'h7456a44b5ed13a7b,64'h53c76871dff702a1,64'hb6f3d259e5fcb53f,
64'h0ea4243a1080115f,64'h62db5c0b9abf8d79,64'he886d57225b6fc7b,64'h8a1ed2c254b2a044,
64'hfafdf655f12048fc,64'h74e90a393ac46233,64'hd8d4b5fe834bb1b1,64'h9f4aafc7a4a6b395,
64'h3affc20312cbe38b,64'h3b0d463d6552a871,64'h83d81879d53d7de7,64'hfffffeff00000101,
64'h11648c88e947c9c0,64'ha159d4aa97656412,64'he133b88f683a2d23,64'he886136f744bd6bc,
64'h117c8eaedf3642c5,64'hace3f76c3b1e55b1,64'h10fb8f115205a66c,64'h7bf05c803ac5c620,
64'hb2573730b9aeeb02,64'h22aca14788021f34,64'h531563ef8bdc494d,64'h379be8bf1e8efb83,
64'h32256fc7aa655c6c,64'hc5420434cbd317b9,64'h30c9343940fb5dd1,64'h40003fffc0000000,
64'h2fb3c4e5e4eec6e9,64'hae8ad488cbda2750,64'hea78ed0d5bfee055,64'h36de7a4b1cbf96a8,
64'h21d484872210022c,64'hec5b6b809357f1b0,64'hbd10daada4b6df90,64'h9143da57ca965409,
64'h9f5fbeca3e240920,64'hae9d214687588c47,64'hfb1a96bef0697637,64'h73e955f89494d673,
64'ha75ff83fc2597c72,64'he761a8c6ccaa550f,64'h307b030f1aa7afbd,64'hffffffdf00000021,
64'h022c91911d28f938,64'hd42b3a9492ecac83,64'hbc2677114d0745a5,64'h9d10c26d6e897ad8,
64'h622f91d57be6c859,64'hf59c7eeca763cab7,64'h821f71e1aa40b4ce,64'h0f7e0b900758b8c4,
64'hd64ae6e55735dd61,64'h84559428710043e7,64'h6a62ac7d917b892a,64'ha6f37d1743d1df71,
64'h8644adf8754cab8e,64'hf8a84085b97a62f8,64'he6192686481f6bbb,64'h080007fff8000000,
64'he5f6789bdc9dd8de,64'h15d15a91197b44ea,64'h7d4f1da14b7fdc0b,64'h06dbcf496397f2d5,
64'h843a909064420046,64'h1d8b6d70126afe36,64'h17a21b55b496dbf2,64'hf2287b4a1952ca82,
64'h13ebf7d947c48124,64'h35d3a428b0eb1189,64'h3f6352d7be0d2ec7,64'hae7d2abe72929acf,
64'hd4ebff07384b2f8f,64'h3cec3518b9954aa2,64'h660f60618354f5f8,64'hfffffffb00000005,
64'h0045923223a51f27,64'hba856751f25d9591,64'h7784cee1c9a0e8b5,64'h13a2184dadd12f5b,
64'hec45f239cf7cd90c,64'h3eb38fdd74ec7957,64'h5043ee3bf548169a,64'h81efc17180eb1719,
64'hfac95cdbcae6bbad,64'h308ab284ee20087d,64'hcd4c558ef22f7126,64'hf4de6fa2087a3bef,
64'h50c895becea99572,64'h1f150810b72f4c5f,64'hbcc324d02903ed78,64'h010000ffff000000,
64'h5cbecf133b93bb1c,64'hc2ba2b51632f689e,64'hafa9e3b3896ffb82,64'h60db79e8cc72fe5b,
64'h50875211cc884009,64'h43b16dadc24d5fc7,64'hc2f44369f692db7f,64'hde450f68832a5951,
64'h827d7efaa8f89025,64'he6ba7484361d6232,64'h27ec6a5ad7c1a5d9,64'h35cfa557ae52535a,
64'h3a9d7fe0c70965f2,64'hc79d86a25732a955,64'h0cc1ec0c306a9ebf,64'h7fffffff00000001,
64'h2008b2462474a3e5,64'hf750ace95e4bb2b3,64'h6ef099dbd9341d17,64'ha274430915ba25ec,
64'h9d88be46b9ef9b22,64'h27d671fb8e9d8f2b,64'hca087dc6bea902d4,64'hf03df82d501d62e4,
64'h7f592b9b195cd776,64'h661156503dc40110,64'h59a98ab19e45ee25,64'h3e9bcdf4210f477e,
64'hca1912b719d532af,64'h23e2a101f6e5e98c,64'h1798649a05207daf,64'h0020001fffe00000,
64'h8b97d9e1e7727764,64'h58574569ec65ed14,64'hd5f53c75b12dff71,64'hac1b6f3c798e5fcc,
64'hea10ea4159910802,64'h28762db59849abf9,64'h385e886d1ed25b70,64'hfbc8a1ec30654b2b,
64'h704fafdef51f1205,64'hdcd74e8fc6c3ac47,64'he4fd8d4a7af834bc,64'hc6b9f4aa35ca4a6c,
64'hc753affb58e12cbf,64'h78f3b0d3eae6552b,64'h21983d81660d53d8,64'hefffffff00000001,
64'h64011648648e947d,64'hbeea159c8bc97657,64'h2dde133b5b2683a3,64'h944e8860a2b744be,
64'hd3b117c8173df365,64'ha4face3ed1d3b1e6,64'h99410fb857d5205b,64'h9e07bf052a03ac5d,
64'h4feb2573232b9aef,64'h0cc22aca07b88022,64'h6b353155d3c8bdc5,64'h47d379be4421e8f0,
64'h39432256c33aa656,64'h847c541fbedcbd32,64'h22f30c9320a40fb6,64'h00040003fffc0000,
64'h9172fb3bbcee4eed,64'h8b0ae8acbd8cbda3,64'hfabea78dd625bfef,64'h95836de70f31cbfa,
64'hdd421d476b322101,64'he50ec5b5d3093580,64'h070bd10da3da4b6e,64'hbf79143ce60ca966,
64'h6e09f5fb7ea3e241,64'h3b9ae9d1d8d87589,64'h9c9fb1a8cf5f0698,64'h98d73e94c6b9494e,
64'h38ea75ff4b1c2598,64'haf1e7619dd5ccaa6,64'h043307b02cc1aa7b,64'hfdffffff00000001,
64'h6c8022c8ac91d290,64'h37dd42b371792ecb,64'ha5bbc266cb64d075,64'h5289d10bd456e898,
64'h7a7622f8a2e7be6d,64'h549f59c79a3a763d,64'hb32821f66afaa40c,64'h73c0f7e04540758c,
64'h29fd64ae4465735e,64'hc198455880f71005,64'h6d66a62a5a7917b9,64'h08fa6f37c8843d1e,
64'h4728644a986754cb,64'hd08f8a8337db97a7,64'h445e6192241481f7,64'h000080007fff8000,
64'h722e5f67179dc9de,64'hb1615d14f7b197b5,64'h3f57d4f19ac4b7fe,64'hd2b06dbc21e63980,
64'hfba843a80d664421,64'h1ca1d8b6ba6126b0,64'h40e17a21747b496e,64'h57ef22875cc1952d,
64'hedc13ebe8fd47c49,64'he7735d395b1b0eb2,64'h1393f63519ebe0d3,64'h531ae7d258d7292a,
64'h071d4ebfe96384b3,64'h55e3cec2fbab9955,64'ha08660f565983550,64'hffbfffff00000001,
64'h0d90045915923a52,64'ha6fba855ce2f25da,64'h74b7784c796c9a0f,64'h0a513a217a8add13,
64'h6f4ec45eb45cf7ce,64'h6a93eb3893474ec8,64'h9665043e4d5f5482,64'h8e781efb88a80eb2,
64'h453fac95888cae6c,64'h783308aab01ee201,64'hedacd4c46b4f22f8,64'h411f4de6b91087a4,
64'ha8e50c88b30cea9a,64'h3a11f15046fb72f5,64'h288bcc322482903f,64'h000010000ffff000,
64'h4e45cbeca2f3b93c,64'h762c2ba23ef632f7,64'h47eafa9df3589700,64'h1a560db7843cc730,
64'hff75087421acc885,64'h03943b16d74c24d6,64'h481c2f43ee8f692e,64'h6afde4508b9832a6,
64'hfdb827d6f1fa8f8a,64'hdcee6ba66b6361d7,64'ha2727ec6033d7c1b,64'hca635cf98b1ae526,
64'ha0e3a9d75d2c7097,64'h6abc79d7ff75732b,64'h1410cc1eacb306aa,64'hfff7ffff00000001,
64'hc1b2008a62b2474b,64'hd4df7509f9c5e4bc,64'h2e96ef096f2d9342,64'ha14a27438f515ba3,
64'h4de9d88b968b9efa,64'h0d527d671268e9d9,64'hd2cca08709abea91,64'hd1cf03deb11501d7,
64'h88a7f592311195ce,64'hef0661147603dc41,64'h1db59a988d69e45f,64'h8823e9bc572210f5,
64'hd51ca19056619d54,64'h67423e29a8df6e5f,64'h2511798624905208,64'h0000020001fffe00,
64'h89c8b97d145e7728,64'h2ec5857427dec65f,64'h08fd5f53be6b12e0,64'h034ac1b6f08798e6,
64'h7feea10e24359911,64'h407287629ae9849b,64'h490385e83dd1ed26,64'h4d5fbc89d1730655,
64'hdfb704fa1e3f51f2,64'h3b9dcd74ad6c6c3b,64'hb44e4fd82067af84,64'h594c6b9ef1635ca5,
64'h341c753acba58e13,64'had578f3a5feeae66,64'hc2821983159660d6,64'hfffeffff00000001,
64'hb8364010ac5648ea,64'h9a9beea0bf38bc98,64'hc5d2dde06de5b269,64'hb42944e7d1ea2b75,
64'hc9bd3b10b2d173e0,64'he1aa4fac024d1d3c,64'hfa59941001357d53,64'h3a39e07bb622a03b,
64'h5114feb2062232ba,64'hfde0cc21aec07b89,64'h23b6b352f1ad3c8c,64'h71047d372ae4421f,
64'h9aa394318acc33ab,64'h2ce847c5151bedcc,64'h04a22f30c4920a41,64'h00000040003fffc0,
64'h1139172fa28bcee5,64'h25d8b0ae64fbd8cc,64'h011fabea77cd625c,64'h406958369e10f31d,
64'heffdd420e486b323,64'ha80e50ebb35d3094,64'h492070bcc7ba3da5,64'h69abf790da2e60cb,
64'hdbf6e09e83c7ea3f,64'ha773b9adf5ad8d88,64'h9689c9fa840cf5f1,64'h6b298d737e2c6b95,
64'ha6838ea6b974b1c3,64'h55aaf1e70bfdd5cd,64'h5850433022b2cc1b,64'hffffdfff00000001,
64'hd706c801558ac91e,64'h13537dd417e71793,64'hf8ba5bbb2dbcb64e,64'h7685289c9a3d456f,
64'h1937a762165a2e7c,64'h9c3549f50049a3a8,64'hbf4b32816026afab,64'ha7473c0ed6c45408,
64'hca229fd580c44658,64'hffbc198355d80f72,64'h8476d669de35a792,64'h2e208fa6c55c8844,
64'hb354728591598676,64'h859d08f822a37dba,64'he09445e538924149,64'h000000080007fff8,
64'h622722e5945179dd,64'h84bb16154c9f7b1a,64'h8023f57ccef9ac4c,64'h680d2b0673c21e64,
64'hbdffba837c90d665,64'h9501ca1cf66ba613,64'h69240e1738f747b5,64'had357ef17b45cc1a,
64'h3b7edc13b078fd48,64'h14ee7735beb5b1b1,64'hf2d1393e70819ebf,64'h6d6531ae0fc58d73,
64'hb4d071d4372e9639,64'h6ab55e3c817fbaba,64'hab0a086564565984,64'hfffffbff00000001,
64'h5ae0d8ffeab15924,64'ha26a6fb9e2fce2f3,64'h5f174b7725b796ca,64'h2ed0a5137347a8ae,
64'h8326f4ebc2cb45d0,64'h1386a93ea0093475,64'hb7e9664f8c04d5f6,64'h14e8e781dad88a81,
64'h194453fab01888cb,64'hdff7832faabb01ef,64'hd08edacc7bc6b4f3,64'h85c411f458ab9109,
64'h566a8e50722b30cf,64'hd0b3a11e44546fb8,64'hfc1288bbc712482a,64'h000000010000ffff,
64'h6c44e45c528a2f3c,64'hd09762c1e993ef64,64'h90047eaf19df358a,64'h8d01a5604e7843cd,
64'h77bff7500f921acd,64'hb2a03942fecd74c3,64'h6d2481c2871ee8f7,64'hd5a6afdd6f68b984,
64'h076fdb82760f1fa9,64'he29dcee5d7d6b637,64'h3e5a2727ae1033d8,64'hadaca63521f8b1af,
64'hf69a0e39a6e5d2c8,64'hcd56abc6d02ff758,64'h9561410c2c8acb31,64'hffffff7f00000001,
64'h8b5c1b1f7d562b25,64'hb44d4df69c5f9c5f,64'hcbe2e96e24b6f2da,64'h45da14a22e68f516,
64'h1064de9d785968ba,64'h6270d5277401268f,64'h56fd2cc9b1809abf,64'he29d1cef5b5b1151,
64'ha3288a7eb603111a,64'h3bfef065d557603e,64'hba11db58ef78d69f,64'hf0b8823dab157222,
64'h2acd51c9ee45661a,64'h1a167423c88a8df7,64'hdf825116b8e24906,64'h2000000000002000,
64'h8d889c8b0a5145e8,64'h9a12ec57bd327ded,64'hd2008fd5233be6b2,64'h71a034aba9cf087a,
64'h6ef7fee9a1f2435a,64'hb6540727bfd9ae99,64'h2da4903830e3dd1f,64'h9ab4d5fb2ded1731,
64'he0edfb6f6ec1e3f6,64'h3c53b9dc9afad6c7,64'h07cb44e4f5c2067b,64'h35b594c6843f1636,
64'h1ed341c734dcba59,64'h19aad578da05feeb,64'hf2ac2820a5915967,64'hffffffef00000001,
64'h716b83638faac565,64'h3689a9beb38bf38c,64'hd97c5d2d0496de5c,64'h48bb429405cd1ea3,
64'hc20c9bd2ef0b2d18,64'h2c4e1aa4ce8024d2,64'h2adfa59916301358,64'hfc53a39d0b6b622b,
64'hd465114f16c06224,64'h477fde0c7aaaec08,64'h37423b6afdef1ad4,64'hde171046f562ae45,
64'hc559aa387dc8acc4,64'h2342ce84591151bf,64'h5bf04a22971c4921,64'h0400000000000400,
64'h11b11391614a28bd,64'h73425d8a97a64fbe,64'hda4011f9e4677cd7,64'hce340694b539e110,
64'hcddeffdc743e486c,64'hf6ca80e417fb35d4,64'h25b49206e61c7ba4,64'hf3569abe85bda2e7,
64'h5c1dbf6dadd83c7f,64'h278a773b735f5ad9,64'ha0f9689bfeb840d0,64'h46b6b2989087e2c7,
64'he3da6838069b974c,64'ha3355aae7b40bfde,64'h3e558503f4b22b2d,64'hfffffffd00000001,
64'h6e2d706c11f558ad,64'h86d1353756717e72,64'h9b2f8ba52092dbcc,64'ha9176851e0b9a3d5,
64'h1841937a5de165a3,64'hc589c353d9d0049b,64'h055bf4b322c6026b,64'hbf8a7473016d6c46,
64'h9a8ca22962d80c45,64'h08effbc18f555d81,64'h86e8476cdfbde35b,64'h7bc2e2087eac55c9,
64'h98ab35468fb91599,64'h246859d06b222a38,64'heb7e094372e38925,64'h0080000000000080,
64'h62362271cc294518,64'h4e684bb112f4c9f8,64'h3b48023f1c8cef9b,64'h19c680d296a73c22,
64'h99bbdffb0e87c90e,64'h9ed9501c02ff66bb,64'h84b692405cc38f75,64'h3e6ad357b0b7b45d,
64'h2b83b7ed95bb0790,64'he4f14ee68e6beb5c,64'h141f2d137fd7081a,64'h28d6d652f210fc59,
64'h9c7b4d0680d372ea,64'h5466ab558f6817fc,64'h67cab0a01e964566,64'hfffffffec0000001,
64'h6dc5ae0d223eab16,64'hd0da26a62ace2fcf,64'h9365f17424125b7a,64'h7522ed09dc17347b,
64'ha308326eabbc2cb5,64'hb8b13869db3a0094,64'ha0ab7e95c458c04e,64'h57f14e8e202dad89,
64'h73519444cc5b0189,64'he11dff7751eaabb1,64'hb0dd08ecfbf7bc6c,64'hef785c402fd58aba,
64'hf31566a7f1f722b4,64'h048d0b3a0d644547,64'h7d6fc1280e5c7125,64'h0010000000000010,
64'h0c46c44e398528a3,64'h09cd0976225e993f,64'ha769004743919df4,64'hc338d01992d4e785,
64'h53377bff21d0f922,64'hb3db2a02e05fecd8,64'h7096d247ab9871ef,64'h67cd5a6a9616f68c,
64'h057076fdb2b760f2,64'h9c9e29dc51cd7d6c,64'hc283e5a1affae104,64'he51adac97e421f8c,
64'hd38f69a0101a6e5e,64'h8a8cd56a31ed0300,64'h4cf95613c3d2c8ad,64'hfffffffef8000001,
64'h4db8b5c16447d563,64'h3a1b44d4a559c5fa,64'hd26cbe2dc4824b70,64'haea45da09b82e690,
64'h7461064d75778597,64'h9716270cbb674013,64'h54156fd2788b180a,64'heafe29d0e405b5b2,
64'hee6a3287b98b6032,64'hfc23bfee0a3d5577,64'h961ba11d1f7ef78e,64'hddef0b8745fab158,
64'h9e62acd47e3ee457,64'h2091a16721ac88a9,64'h6fadf824a1cb8e25,64'h0002000000000002,
64'ha188d8892730a515,64'h2139a12ea44bd328,64'h94ed2008687233bf,64'h78671a02d25a9cf1,
64'hca66ef7f243a1f25,64'h167b65405c0bfd9b,64'h2e12da48d5730e3e,64'h8cf9ab4cd2c2ded2,
64'hc0ae0edef656ec1f,64'h9393c53b0a39afae,64'h98507cb3b5ff5c21,64'h9ca35b58afc843f2,
64'h5a71ed33c2034dcc,64'h11519aad463da060,64'h699f2ac2187a5916,64'hfffffffeff000001,
64'ha9b716b78c88faad,64'hc7436899d4ab38c0,64'h1a4d97c5b890496e,64'h15d48bb413705cd2,
64'h2e8c20c98eaef0b3,64'hb2e2c4e0f76ce803,64'hca82adf98f116302,64'hdd5fc5395c80b6b7,
64'hddcd465037316c07,64'h3f8477fda147aaaf,64'h52c3742363efdef2,64'h1bbde170e8bf562b,
64'h33cc559a6fc7dc8b,64'he412342c04359116,64'h6df5bf04343971c5,64'hc0003fff40000001,
64'h74311b10c4e614a3,64'h04273425d4897a65,64'h329da400ed0e4678,64'hef0ce33f7a4b539f,
64'h794cddef848743e5,64'ha2cf6ca76b817fb4,64'h45c25b48daae61c8,64'hd19f3568da585bdb,
64'h3815c1dbbecadd84,64'h527278a7214735f6,64'hf30a0f9596bfeb85,64'hd3946b6a55f9087f,
64'h8b4e3da5f84069ba,64'h022a3355a8c7b40c,64'h4d33e558030f4b23,64'hfffffffeffe00001,
64'h7536e2d691911f56,64'h18e86d133a956718,64'h4349b2f87712092e,64'hc2ba9175c26e0b9b,
64'ha5d1841891d5de17,64'hb65c589b7eed9d01,64'hd95055be71e22c61,64'h3babf8a70b9016d7,
64'h3bb9a8c9e6e62d81,64'h27f08eff9428f556,64'hca586e83ac7dfbdf,64'ha377bc2d7d17eac6,
64'ha6798ab2adf8fb92,64'h5c8246854086b223,64'h6dbeb7e026872e39,64'hf80007ff08000001,
64'hae862361789cc295,64'h6084e6845a912f4d,64'h0653b4801da1c8cf,64'h3de19c67cf496a74,
64'h6f299bbd9090e87d,64'h9459ed946d702ff7,64'h08b84b691b55cc39,64'hba33e6ac7b4b0b7c,
64'h8702b83af7d95bb1,64'h4a4e4f14a428e6bf,64'h7e6141f252d7fd71,64'h3a728d6d2abf2110,
64'hd169c7b3ff080d38,64'h8045466a3518f682,64'ha9a67caa6061e965,64'hfffffffefffc0001,
64'h4ea6dc5a923223eb,64'h031d0da26752ace3,64'h4869365ecee24126,64'hb857522e184dc174,
64'h34ba3082f23abbc3,64'hf6cb8b128fddb3a1,64'hfb2a0ab6ee3c458d,64'h27757f14c17202db,
64'he77735185cdcc5b1,64'h44fe11dfb2851eab,64'h394b0dd0558fbf7c,64'h546ef7856fa2fd59,
64'hd4cf315595bf1f73,64'hab9048d00810d645,64'hedb7d6fb24d0e5c8,64'hff0000ff01000001,
64'h75d0c46bcf139853,64'h6c109cd02b5225ea,64'h20ca768fe3b4391a,64'h87bc338c79e92d4f,
64'h6de5337752121d10,64'h328b3db26dae05ff,64'he117096c436ab988,64'h97467cd50f696170,
64'hf0e057067efb2b77,64'h2949c9e274851cd8,64'hefcc283d6a5affaf,64'h074e51ada557e422,
64'h1a2d38f67fe101a7,64'hd008a8cc86a31ed1,64'h7534cf94ec0c3d2d,64'hfffffffeffff8001,
64'ha9d4db8ab246447e,64'ha063a1b3acea559d,64'h490d26cb99dc4825,64'h970aea454309b82f,
64'ha697460fbe475779,64'hfed9716171fbb675,64'h7f6541567dc788b2,64'ha4eeafe1f82e405c,
64'hfceee6a22b9b98b7,64'ha89fc23b5650a3d6,64'h872961b98ab1f7f0,64'hea8ddeefcdf45fac,
64'hba99e62a12b7e3ef,64'h75720919a1021ac9,64'h1db6fadf649a1cb9,64'hffe0001f00200001,
64'haeba188cd9e2730b,64'hcd821399456a44be,64'hc4194ed13c768724,64'h30f786716f3d25aa,
64'h0dbca66eea4243a2,64'h265167b62db5c0c0,64'h1c22e12d886d5731,64'h12e8cf9aa1ed2c2e,
64'h3e1c0ae0afdf656f,64'h0529393c4e90a39b,64'h3df985078d4b5ff6,64'hc0e9ca34f4aafc85,
64'h2345a71eaffc2035,64'hfa011518b0d463db,64'h6ea699f23d8187a6,64'hfffffffefffff001,
64'h553a9b711648c890,64'h740c7436159d4ab4,64'h6921a4d9133b8905,64'h32e15d4888613706,
64'hf4d2e8c117c8eaf0,64'h7fdb2e2bce3f76cf,64'hcfeca82a0fb8f117,64'h949dd5fbbf05c80c,
64'h3f9ddcd425737317,64'h5513f8472aca147b,64'h10e52c3731563efe,64'h9d51bbdd79be8bf6,
64'h37533cc52256fc7e,64'heeae41225420435a,64'he3b6df5b0c934398,64'hfffc000300040001,
64'hb5d74310fb3c4e62,64'h59b04272e8ad4898,64'h988329d9a78ed0e5,64'hc61ef0cd6de7a4b6,
64'hc1b794cd1d484875,64'h04ca2cf6c5b6b818,64'he3845c24d10daae7,64'h425d19f3143da586,
64'h27c3815bf5fbecae,64'ha0a52726e9d21474,64'h47bf30a0b1a96bff,64'h781d39463e955f91,
64'h6468b4e375ff8407,64'hbf4022a2761a8c7c,64'h4dd4d33e07b030f5,64'hfffffffefffffe01,
64'h0aa7536e22c91912,64'h8e818e8642b3a957,64'h6d24349ac2677121,64'h465c2ba8d10c26e1,
64'h1e9a5d1822f91d5e,64'h2ffb65c559c7eeda,64'h39fd950521f71e23,64'h9293babef7e0b902,
64'h27f3bb9a64ae6e63,64'haaa27f0845594290,64'h421ca586a62ac7e0,64'h53aa377b6f37d17f,
64'h46ea6798644adf90,64'hddd5c8238a84086c,64'h1c76dbeb61926873,64'hffff7fff80008001,
64'hd6bae8615f6789cd,64'h0b36084e5d15a913,64'h7310653ad4f1da1d,64'h58c3de196dbcf497,
64'h7836f29943a9090f,64'h0099459ed8b6d703,64'h3c708b847a21b55d,64'h484ba33e2287b4b1,
64'h44f8702b3ebf7d96,64'h9414a4e45d3a428f,64'h28f7e613f6352d80,64'hef03a727e7d2abf3,
64'h2c8d169c4ebff081,64'h97e80453cec35190,64'h69ba9a6760f6061f,64'hfffffffeffffffc1,
64'hc154ea6d04592323,64'h31d031d0a856752b,64'heda48692784cee25,64'he8cb85743a2184dd,
64'h43d34ba2c45f23ac,64'hc5ff6cb7eb38fddc,64'ha73fb2a0043ee3c5,64'hd25277571efc1721,
64'ha4fe7772ac95cdcd,64'h15544fe108ab2852,64'h084394b0d4c558fc,64'h2a7546ef4de6fa30,
64'h08dd4cf30c895bf2,64'h9bbab903f150810e,64'ha38edb7ccc324d0f,64'hffffefff10001001,
64'h7ad75d0bcbecf13a,64'ha166c1092ba2b523,64'h6e620ca6fa9e3b44,64'h2b187bc30db79e93,
64'h2f06de5308752122,64'ha01328b33b16dae1,64'h678e11702f4436ac,64'he9097466e450f697,
64'h489f0e0527d7efb3,64'h3282949c6ba74852,64'h051efcc27ec6a5b0,64'hbde074e45cfa557f,
64'he591a2d2a9d7fe11,64'h12fd008a79d86a32,64'h2d37534ccc1ec0c4,64'hfffffffefffffff9,
64'hb82a9d4d008b2465,64'ha63a0639750acea6,64'h7db490d1ef099dc5,64'h7d1970ae2744309c,
64'h887a6973d88be476,64'h98bfed967d671fbc,64'h74e7f653a087dc79,64'hfa4a4eea03df82e5,
64'h749fceedf592b9ba,64'hc2aa89fb6115650b,64'h810872959a98ab20,64'h054ea8dde9bcdf46,
64'hc11ba99da1912b7f,64'h537757203e2a1022,64'h3471db6f798649a2,64'hfffffdff02000201,
64'hcf5aeba0b97d9e28,64'hb42cd820857456a5,64'h8dcc41945f53c769,64'ha5630f77c1b6f3d3,
64'hc5e0dbc9a10ea425,64'hf40265158762db5d,64'h8cf1c22d85e886d6,64'h3d212e8cbc8a1ed3,
64'ha913e1c004fafdf7,64'hc6505292cd74e90b,64'h00a3df984fd8d4b6,64'h37bc0e9c6b9f4ab0,
64'hfcb23459753affc3,64'hc25fa0108f3b0d47,64'h85a6ea691983d819,64'hffffffff00000000,
64'h770553a94011648d,64'h54c740c6eea159d5,64'h6fb69219dde133b9,64'h8fa32e1544e88614,
64'h510f4d2e3b117c8f,64'h9317fdb24face3f8,64'hee9cfec99410fb90,64'h7f4949dce07bf05d,
64'hce93f9dcfeb25738,64'hb855513ecc22aca2,64'h10210e52b3531564,64'h40a9d51b7d379be9,
64'h3823753394322570,64'hca6eeae347c54205,64'hc68e3b6d2f30c935,64'hffffffbf00400041,
64'h19eb5d74172fb3c5,64'h76859b03b0ae8ad5,64'hf1b98831abea78ee,64'hb4ac61ee5836de7b,
64'h78bc1b78d421d485,64'h7e804ca250ec5b6c,64'h519e384570bd10db,64'ha7a425d0f79143db,
64'h35227c37e09f5fbf,64'hb8ca0a51b9ae9d22,64'h40147bf2c9fb1a97,64'h06f781d38d73e956,
64'hbf96468a8ea75ff9,64'h384bf401f1e761a9,64'hf0b4dd4c43307b04,64'h1fffffffe0000000,
64'h6ee0aa74c8022c92,64'h6a98e8187dd42b3b,64'hedf6d2425bbc2678,64'h91f465c2289d10c3,
64'h2a21e9a5a7622f92,64'h1262ffb649f59c7f,64'h1dd39fd932821f72,64'h6fe9293b3c0f7e0c,
64'h19d27f3b9fd64ae7,64'hd70aaa2719845595,64'h820421c9d66a62ad,64'he8153aa28fa6f37e,
64'h07046ea6728644ae,64'h794ddd5c08f8a841,64'h78d1c76d45e61927,64'hfffffff700080009,
64'h633d6bae22e5f679,64'h6ed0b3601615d15b,64'h5e373105f57d4f1e,64'hb6958c3d2b06dbd0,
64'h6f17836eba843a91,64'h8fd00993ca1d8b6e,64'haa33c7080e17a21c,64'hb4f484b97ef2287c,
64'h26a44f86dc13ebf8,64'hd71941497735d3a5,64'h28028f7e393f6353,64'h40def03a31ae7d2b,
64'hf7f2c8d071d4ec00,64'he7097e7f5e3cec36,64'h9e169ba908660f61,64'h03fffffffc000000,
64'hcddc154dd9004593,64'had531d026fba8568,64'h1dbeda484b7784cf,64'hb23e8cb7a513a219,
64'hc5443d33f4ec45f3,64'h224c5ff6a93eb390,64'hc3ba73fa665043ef,64'h8dfd2526e781efc2,
64'h233a4fe753fac95d,64'h7ae1554483308ab3,64'h70408438dacd4c56,64'h5d02a75411f4de70,
64'h40e08dd48e50c896,64'hef29bbaaa11f1509,64'h2f1a38ed88bcc325,64'hfffffffe00010002,
64'hec67ad74e45cbed0,64'hadda166b62c2ba2c,64'h4bc6e6207eafa9e4,64'h16d2b187a560db7a,
64'hede2f06cf7508753,64'h51fa01323943b16e,64'h954678e081c2f444,64'h969e9096afde4510,
64'h04d489f0db827d7f,64'h7ae32828cee6ba75,64'ha50051ef2727ec6b,64'ha81bde06a635cfa6,
64'h1efe591a0e3a9d80,64'h5ce12fcfabc79d87,64'hf3c2d374410cc1ed,64'h007fffffff800000,
64'hb9bb82a91b2008b3,64'h15aa63a04df750ad,64'h23b7db48e96ef09a,64'hf647d19614a27444,
64'hb8a887a5de9d88bf,64'h04498bfed527d672,64'h38774e7f2cca087e,64'hd1bfa4a41cf03df9,
64'h646749fc8a7f592c,64'haf5c2aa7f0661157,64'h4e081086db59a98b,64'h0ba054ea823e9bce,
64'h481c11ba51ca1913,64'hfde537747423e2a2,64'h65e3471d51179865,64'hdfffffff00002001,
64'h1d8cf5ae9c8b97da,64'h95bb42ccec585746,64'h8978dcc38fd5f53d,64'hc2da563034ac1b70,
64'hbdbc5e0cfeea10eb,64'h4a3f40260728762e,64'h92a8cf1b90385e89,64'h12d3d212d5fbc8a2,
64'h209a913dfb704fb0,64'h6f5c6504b9dcd74f,64'hb4a00a3d44e4fd8e,64'h55037bc094c6b9f5,
64'h03dfcb2341c753b0,64'h2b9c25f9d578f3b1,64'h7e785a6e2821983e,64'h000ffffffff00000,
64'hb737705483640117,64'h62b54c73a9beea16,64'hc476fb685d2dde14,64'h9ec8fa3242944e89,
64'h371510f49bd3b118,64'hc089317f1aa4facf,64'h470ee9cfa5994110,64'hfa37f493a39e07c0,
64'h8c8ce93f114feb26,64'h35eb8554de0cc22b,64'ha9c102103b6b3532,64'h41740a9d1047d37a,
64'ha9038236aa394323,64'hdfbca6edce847c55,64'h6cbc68e34a22f30d,64'hfbffffff00000401,
64'hc3b19eb5139172fc,64'h52b768595d8b0ae9,64'h712f1b9811fabea8,64'h185b4ac60695836e,
64'hb7b78bc0ffdd421e,64'h4947e80480e50ec6,64'hf25519e292070bd2,64'hc25a7a419abf7915,
64'h04135227bf6e09f6,64'h2deb8ca0773b9aea,64'h56940147689c9fb2,64'h6aa06f77b298d73f,
64'h007bf9646838ea76,64'he57384be5aaf1e77,64'h4fcf0b4d85043308,64'h0001fffffffe0000,
64'h36e6ee0a706c8023,64'h4c56a98e3537dd43,64'h988edf6c8ba5bbc3,64'hf3d91f45685289d2,
64'h06e2a21e937a7623,64'h3811262fc3549f5a,64'h08e1dd39f4b32822,64'h1f46fe927473c0f8,
64'h51919d27a229fd65,64'ha6bd70a9fbc19846,64'hd5382041476d66a7,64'hc82e8152e208fa70,
64'hb520704635472865,64'h7bf794dd59d08f8b,64'h6d978d1c09445e62,64'hff7fffff00000081,
64'h987633d622722e60,64'hea56ed0a4bb1615e,64'h0e25e373023f57d5,64'h430b695880d2b06e,
64'h56f6f177dffba844,64'h4928fd00501ca1d9,64'hde4aa33b9240e17b,64'h784b4f47d357ef23,
64'h40826a44b7edc13f,64'hc5bd71934ee7735e,64'hcad280282d1393f7,64'h2d540deed6531ae8,
64'h400f7f2c4d071d4f,64'h3cae7097ab55e3cf,64'h09f9e169b0a08661,64'h00003fffffffc000,
64'ha6dcddc0ae0d9005,64'ha98ad53126a6fba9,64'hb311dbecf174b779,64'hde7b23e7ed0a513b,
64'ha0dc5443326f4ec5,64'hc70224c5386a93ec,64'hc11c3ba67e966505,64'h03e8dfd24e8e781f,
64'h6a3233a494453fad,64'h54d7ae14ff783309,64'h3aa7040808edacd5,64'h1905d02a5c411f4e,
64'h76a40e0866a8e50d,64'haf7ef29b0b3a11f2,64'hcdb2f1a2c1288bcd,64'hffefffff00000011,
64'h130ec67ac44e45cc,64'h5d4adda109762c2c,64'h61c4bc6e0047eafb,64'h48616d2ad01a560e,
64'h8adede2e7bff7509,64'he9251f9f2a03943c,64'hbbc95466d2481c30,64'haf0969e85a6afde5,
64'h28104d4876fdb828,64'h58b7ae3229dcee6c,64'h395a5004e5a2727f,64'h05aa81bddaca635d,
64'h2801efe569a0e3aa,64'h2795ce12d56abc7a,64'he13f3c2c561410cd,64'h000007fffffff800,
64'h74db9bb7b5c1b201,64'hf5315aa544d4df76,64'hf6623b7cbe2e96f0,64'hbbcf647c5da14a28,
64'h741b8a88064de9d9,64'h98e04498270d527e,64'h782387746fd2cca1,64'h207d1bfa29d1cf04,
64'h6d4646743288a7f6,64'hea9af5c1bfef0662,64'h6754e080a11db59b,64'h4320ba050b8823ea,
64'h6ed481c0acd51ca2,64'hd5efde52a167423f,64'h79b65e33f825117a,64'hfffdffff00000003,
64'h8261d8ced889c8ba,64'h8ba95bb3a12ec586,64'hac38978d2008fd60,64'h490c2da51a034ac2,
64'hf15bdbc4ef7feea2,64'h9d24a3f365407288,64'h17792a8cda490386,64'h75e12d3cab4d5fbd,
64'h050209a90edfb705,64'h8b16f5c5c53b9dce,64'h272b4a007cb44e50,64'h60b550375b594c6c,
64'hc5003dfbed341c76,64'hc4f2b9c19aad5790,64'h7c27e7852ac2821a,64'h000000ffffffff00,
64'hee9b737616b83641,64'h5ea62b54689a9bef,64'h1ecc476f97c5d2de,64'h1779ec8f8bb42945,
64'hee83715020c9bd3c,64'h531c0892c4e1aa50,64'hef0470edadfa5995,64'h840fa37ec53a39e1,
64'h4da8c8ce465114ff,64'hdd535eb777fde0cd,64'hacea9c0f7423b6b4,64'hc864173fe171047e,
64'hcdda9037559aa395,64'h3abdfbca342ce848,64'hcf36cbc5bf04a230,64'hbfffbfff40000001,
64'hd04c3b191b113918,64'h51752b763425d8b1,64'h158712f1a4011fac,64'hc92185b3e3406959,
64'hde2b7b77ddeffdd5,64'h13a4947e6ca80e51,64'h42ef25515b492071,64'h6ebc25a73569abf8,
64'h60a04134c1dbf6e1,64'h5162deb878a773ba,64'h04e569400f9689ca,64'h8c16aa066b6b298e,
64'h58a007bf3da6838f,64'h189e57383355aaf2,64'hcf84fcefe5585044,64'h0000001fffffffe0,
64'hfdd36e6de2d706c9,64'h2bd4c56a6d13537e,64'h43d988edb2f8ba5c,64'h62ef3d9191768529,
64'h9dd06e29841937a8,64'h0a638112589c354a,64'h7de08e1d55bf4b33,64'hf081f46ef8a7473d,
64'h29b51919a8ca22a0,64'h7baa6bd68effbc1a,64'h959d53816e8476d7,64'h590c82e7bc2e2090,
64'h79bb52068ab35473,64'h0757bf7946859d09,64'h19e6d978b7e09446,64'hf7fff7ff08000001,
64'h1a09876323622723,64'hea2ea56de684bb17,64'h82b0e25db48023f6,64'hf92430b59c680d2c,
64'h7bc56f6e9bbdffbb,64'he274928eed9501cb,64'he85de4a94b69240f,64'h0dd784b4e6ad357f,
64'hec140825b83b7edd,64'hca2c5bd64f14ee78,64'hc09cad2741f2d13a,64'h5182d5408d6d6532,
64'h2b1400f7c7b4d072,64'hc313cae6466ab55f,64'h99f09f9d7cab0a09,64'h00000003fffffffc,
64'hffba6dccdc5ae0da,64'h457a98ad0da26a70,64'h887b311d365f174c,64'hec5de7b1522ed0a6,
64'h13ba0dc5308326f5,64'hc14c70218b1386aa,64'hafbc11c30ab7e967,64'h7e103e8d7f14e8e8,
64'h0536a32335194454,64'hcf754d7a11dff784,64'h32b3aa700dd08edb,64'h0b21905cf785c412,
64'haf376a4031566a8f,64'he0eaf7ee48d0b3a2,64'h433cdb2ed6fc1289,64'hfefffeff01000001,
64'ha34130ebc46c44e5,64'h3d45d4ad9cd09763,64'h50561c4b7690047f,64'h9f248616338d01a6,
64'haf78aded3377bff8,64'hbc4e92513db2a03a,64'h3d0bbc95096d2482,64'h21baf0967cd5a6b0,
64'h7d82810457076fdc,64'h19458b7ac9e29dcf,64'hd81395a4283e5a28,64'hca305aa751adaca7,
64'hc562801e38f69a0f,64'h3862795ca8cd56ac,64'hf33e13f2cf956142,64'h8000000000000000,
64'hdff74db8db8b5c1c,64'h08af5315a1b44d4e,64'h910f662326cbe2ea,64'h5d8bbcf5ea45da15,
64'h627741b8461064df,64'hd8298e03716270d6,64'h35f782384156fd2d,64'h0fc207d1afe29d1d,
64'h80a6d463e6a3288b,64'h99eea9aec23bfef1,64'ha656754d61ba11dc,64'hc164320adef0b883,
64'h35e6ed47e62acd52,64'hdc1d5efd091a1675,64'he8679b64fadf8252,64'hffdfffdf00200001,
64'h7468261d188d889d,64'ha7a8ba95139a12ed,64'h2a0ac3894ed20090,64'h53e490c28671a035,
64'h15ef15bda66ef7ff,64'hd789d24967b65408,64'hc7a17791e12da491,64'h04375e12cf9ab4d6,
64'h8fb050200ae0edfc,64'h2328b16f393c53ba,64'h1b0272b48507cb45,64'h39460b54ca35b595,
64'h38ac5003a71ed342,64'h870c4f2b1519aad6,64'hde67c27d99f2ac29,64'h1000000000000000,
64'h9bfee9b69b716b84,64'h4115ea62743689aa,64'hd221ecc3a4d97c5e,64'h6bb1779e5d48bb43,
64'h2c4ee836e8c20c9c,64'h5b0531c02e2c4e1b,64'h66bef046a82adfa6,64'h61f840f9d5fc53a4,
64'hb014da8bdcd46512,64'hf33dd534f8477fdf,64'h94cacea92c37423c,64'hb82c8640bbde1711,
64'hc6bcdda83cc559ab,64'h7b83abdf412342cf,64'hdd0cf36bdf5bf04b,64'hfffbfffb00040001,
64'h6e8d04c34311b114,64'h74f517524273425e,64'h0541587129da4012,64'h6a7c9217f0ce3407,
64'h22bde2b794cddf00,64'h1af13a492cf6ca81,64'hf8f42ef15c25b493,64'h4086ebc219f3569b,
64'h91f60a03815c1dc0,64'hc465162d27278a78,64'h63604e5630a0f969,64'h6728c16a3946b6b3,
64'hc71589ffb4e3da69,64'h50e189e522a3355b,64'hfbccf84ed33e5586,64'h0200000000000000,
64'h937fdd36536e2d71,64'hc822bd4b8e86d136,64'h5a443d98349b2f8c,64'had762ef32ba91769,
64'h8589dd065d184194,64'hab60a63765c589c4,64'h4cd7de0895055bf5,64'h8c3f081ebabf8a75,
64'hd6029b50bb9a8ca3,64'h3e67baa67f08effc,64'h929959d4a586e848,64'hf70590c7377bc2e3,
64'hb8d79bb46798ab36,64'h2f70757bc824685a,64'hbba19e6cdbeb7e0a,64'hffff7ffe80008001,
64'h8dd1a097e8623623,64'h4e9ea2ea084e684c,64'hc0a82b0d653b4803,64'h2d4f9242de19c681,
64'h0457bc56f299bbe0,64'he35e2748459ed951,64'hbf1e85dd8b84b693,64'ha810dd77a33e6ad4,
64'h123ec140702b83b8,64'h188ca2c5a4e4f14f,64'hec6c09c9e6141f2e,64'hace5182ca728d6d7,
64'hf8e2b13f169c7b4e,64'haa1c313c045466ac,64'h5f799f099a67cab1,64'h0040000000000000,
64'hf26ffba5ea6dc5af,64'h590457a931d0da27,64'h8b4887b2869365f2,64'hf5aec5dd857522ee,
64'h90b13ba04ba30833,64'h956c14c66cb8b139,64'h699afbc0b2a0ab7f,64'h7187e1037757f14f,
64'hbac0536977735195,64'h87ccf7544fe11e00,64'h12532b3a94b0dd09,64'hbee0b21846ef785d,
64'h571af3764cf31567,64'hc5ee0eaeb9048d0c,64'hd77433ccdb7d6fc2,64'hffffeffef0001001,
64'hb1ba34125d0c46c5,64'h89d3d45cc109cd0a,64'hb81505610ca76901,64'he5a9f2477bc338d1,
64'h008af78ade53377c,64'hfc6bc4e828b3db2b,64'hb7e3d0bb117096d3,64'h95021bae7467cd5b,
64'h0247d8280e057077,64'h23119458949c9e2a,64'h5d8d8138fcc283e6,64'h359ca30574e51adb,
64'h5f1c5627a2d38f6a,64'h95438627008a8cd6,64'hebef33e0534cf957,64'h0008000000000000,
64'h3e4dff749d4db8b6,64'h2b208af5063a1b45,64'hd16910f590d26cbf,64'h5eb5d8bb70aea45e,
64'hb216277369746107,64'hf2ad8297ed971628,64'h2d335f77f6541570,64'h2e30fc204eeafe2a,
64'h77580a6cceee6a33,64'h10f99eea89fc23c0,64'he24a656672961ba2,64'h77dc1642a8ddef0c,
64'h2ae35e6ea99e62ad,64'h98bdc1d5572091a2,64'hdaee8678db6fadf9,64'hfffffdfefe000201,
64'h76374681eba188d9,64'hd13a7a8ad82139a2,64'hf702a0ab4194ed21,64'hfcb53e480f78671b,
64'h80115ef0dbca66f0,64'hbf8d789c65167b66,64'hb6fc7a16c22e12db,64'hb2a043752e8cf9ac,
64'h2048fb04e1c0ae0f,64'hc462328a529393c6,64'h4bb1b026df98507d,64'ha6b394600e9ca35c,
64'hcbe38ac4345a71ee,64'h52a870c4a011519b,64'h3d7de67bea699f2b,64'h0001000000000000,
64'h47c9bfee53a9b717,64'h6564115e40c74369,64'h3a2d221e921a4d98,64'h4bd6bb172e15d48c,
64'h3642c4ee4d2e8c21,64'h1e55b052fdb2e2c5,64'h05a66beefeca82ae,64'hc5c61f8349dd5fc6,
64'haeeb014cf9ddcd47,64'h021f33dd513f8478,64'hdc494cac0e52c375,64'h8efb82c7d51bbde2,
64'h655c6bcd7533cc56,64'hd317b839eae41235,64'hfb5dd0ce3b6df5c0,64'hffffffbeffc00041,
64'heec6e8cf5d74311c,64'hda274f509b042735,64'hfee0541488329da5,64'hbf96a7c861ef0ce4,
64'h10022bde1b794cde,64'h57f1af134ca2cf6d,64'hb6df8f423845c25c,64'h9654086e25d19f36,
64'h24091f607c3815c2,64'h588c46510a527279,64'h697636047bf30a10,64'h94d6728b81d3946c,
64'h597c7158468b4e3e,64'haa550e17f4022a34,64'ha7afbccedd4d33e6,64'h0000200000000000,
64'h28f937fdaa7536e3,64'hecac822ae818e86e,64'h0745a443d24349b3,64'h897ad76265c2ba92,
64'he6c8589ce9a5d185,64'h63cab609ffb65c59,64'h40b4cd7d9fd95056,64'h58b8c3f0293babf9,
64'h35dd60297f3bb9a9,64'h0043e67baa27f08f,64'h7b89299521ca586f,64'hd1df70583aa377bd,
64'h4cab8d796ea6798b,64'h7a62f706dd5c8247,64'h1f6bba19c76dbeb8,64'hfffffff6fff80009,
64'h9dd8dd196bae8624,64'h7b44e9e9b36084e7,64'h7fdc0a82310653b5,64'h97f2d4f88c3de19d,
64'h4200457b836f299c,64'h6afe35e2099459ee,64'h96dbf1e7c708b84c,64'h52ca810d84ba33e7,
64'hc48123eb4f8702b9,64'heb1188c9414a4e50,64'h0d2ec6c08f7e6142,64'h929ace50f03a728e,
64'h4b2f8e2ac8d169c8,64'h954aa1c27e804547,64'h54f5f7999ba9a67d,64'h0000040000000000,
64'ha51f26ff154ea6dd,64'h5d9590451d031d0e,64'ha0e8b487da486937,64'hd12f5aeb8cb85753,
64'h7cd90b133d34ba31,64'hec7956c05ff6cb8c,64'h481699af73fb2a0b,64'heb17187d25277580,
64'he6bbac044fe77736,64'h20087ccf5544fe12,64'h2f71253284394b0e,64'h7a3bee0aa7546ef8,
64'ha99571ae8dd4cf32,64'h2f4c5ee0bbab9049,64'h03ed774338edb7d7,64'hfffffffdffff0002,
64'h93bb1ba2ad75d0c5,64'h2f689d3d166c109d,64'h6ffb814fe620ca77,64'h72fe5a9eb187bc34,
64'h884008aef06de534,64'h4d5fc6bc01328b3e,64'h92db7e3c78e1170a,64'h2a5950219097467d,
64'hf890247c89f0e058,64'h1d623119282949ca,64'hc1a5d8d751efcc29,64'h525359c9de074e52,
64'h0965f1c5591a2d39,64'h32a954382fd008a9,64'h6a9ebef2d37534d0,64'h0000008000000000,
64'h74a3e4df82a9d4dc,64'h4bb2b20863a063a2,64'h341d1690db490d27,64'hba25eb5cd1970aeb,
64'hef9b216187a69747,64'h9d8f2ad78bfed972,64'ha902d3354e7f6542,64'h1d62e30fa4a4eeb0,
64'h5cd7758049fceee7,64'hc4010f992aa89fc3,64'h45ee24a610872962,64'h0f477dc154ea8ddf,
64'hd532ae3511ba99e7,64'he5e98bdb3775720a,64'h207daee8471db6fb,64'hdffffffeffffe001,
64'h72776373f5aeba19,64'h65ed13a742cd8214,64'h2dff7029dcc4194f,64'h8e5fcb535630f787,
64'h910801155e0dbca7,64'h49abf8d740265168,64'hd25b6fc6cf1c22e2,64'h654b2a03d212e8d0,
64'h1f12048f913e1c0b,64'hc3ac46226505293a,64'hf834bb1a0a3df986,64'hca4a6b387bc0e9cb,
64'he12cbe37cb2345a8,64'he6552a8625fa0116,64'h0d53d7de5a6ea69a,64'h0000001000000000,
64'h8e947c9b70553a9c,64'hc97656404c740c75,64'h2683a2d1fb6921a5,64'hb744bd6afa32e15e,
64'h3df3642c10f4d2e9,64'hd3b1e55a317fdb2f,64'hd5205a65e9cfeca9,64'h03ac5c61f4949dd6,
64'h2b9aeeafe93f9ddd,64'hb88021f2855513f9,64'hc8bdc4940210e52d,64'h21e8efb80a9d51bc,
64'h3aa655c68237533d,64'hdcbd317aa6eeae42,64'ha40fb5dc68e3b6e0,64'hfbfffffefffffc01,
64'hee4eec6d9eb5d744,64'h8cbda2746859b043,64'h25bfee051b98832a,64'h31cbf96a4ac61ef1,
64'h322100228bc1b795,64'h09357f1ae804ca2d,64'hda4b6df819e3845d,64'h0ca965407a425d1a,
64'ha3e240915227c382,64'hd87588c38ca0a528,64'h5f0697630147bf31,64'hb9494d666f781d3a,
64'h1c2597c6f96468b5,64'h5ccaa55084bf4023,64'hc1aa7afb0b4dd4d4,64'h0000000200000000,
64'h91d28f92ee0aa754,64'h792ecac7a98e818f,64'h64d07459df6d2435,64'h56e897ad1f465c2c,
64'he7be6c84a21e9a5e,64'h3a763cab262ffb66,64'hfaa40b4bdd39fd96,64'h40758b8bfe9293bb,
64'h65735dd59d27f3bc,64'hf710043d70aaa280,64'h7917b89220421ca6,64'h843d1df68153aa38,
64'h6754cab87046ea68,64'hdb97a62e94ddd5c9,64'h1481f6bb8d1c76dc,64'hff7ffffeffffff81,
64'h9dc9dd8d33d6bae9,64'hb197b44ded0b3609,64'hc4b7fdbfe3731066,64'he6397f2c6958c3df,
64'h66442003f17836f3,64'h6126afe2fd009946,64'h7b496dbea33c708c,64'hc1952ca74f484ba4,
64'hd47c48116a44f871,64'h1b0eb118719414a5,64'hebe0d2eb8028f7e7,64'hd72929ac0def03a8,
64'h6384b2f87f2c8d17,64'hab9954a97097e805,64'h98354f5ee169ba9b,64'h0000000040000000,
64'h923a51f1ddc154eb,64'h2f25d958d531d032,64'h6c9a0e8adbeda487,64'h8add12f523e8cb86,
64'h5cf7cd905443d34c,64'h474ec79524c5ff6d,64'h5f5481693ba73fb3,64'ha80eb170dfd25278,
64'h8cae6bba33a4fe78,64'h1ee20087ae155450,64'h4f22f71204084395,64'h1087a3bed02a7547,
64'h0cea99570e08dd4d,64'hfb72f4c4f29bbaba,64'h82903ed6f1a38edc,64'hffeffffefffffff1,
64'hf3b93bb0c67ad75e,64'hf632f688dda166c2,64'h5896ffb7bc6e620d,64'h3cc72fe56d2b187c,
64'hacc883ffde2f06df,64'h4c24d5fc1fa01329,64'h8f692db754678e12,64'h9832a59469e90975,
64'hfa8f89014d489f0f,64'h6361d622ae328295,64'h3d7c1a5d50051efd,64'h1ae5253581bde075,
64'h2c70965eefe591a3,64'h75732a94ce12fd01,64'hb306a9eb3c2d3754,64'h0000000008000000,
64'hb2474a3d9bb82a9e,64'hc5e4bb2a5aa63a07,64'h2d9341d13b7db491,64'h515ba25e647d1971,
64'h8b9ef9b18a887a6a,64'h68e9d8f24498bfee,64'habea902c8774e7f7,64'h1501d62e1bfa4a4f,
64'h1195cd7746749fcf,64'h03dc4010f5c2aa8a,64'h69e45ee1e0810873,64'h2210f477ba054ea9,
64'h619d532a81c11baa,64'hdf6e5e97de537758,64'h905207da5e3471dc,64'hfffdfffeffffffff,
64'h5e772775d8cf5aec,64'hdec65ed05bb42cd9,64'h6b12dff6978dcc42,64'h8798e5fc2da56310,
64'h3599107fdbc5e0dc,64'he9849abea3f40266,64'hd1ed25b62a8cf1c3,64'h730654b22d3d212f,
64'h3f51f12009a913e2,64'h6c6c3ac3f5c65053,64'h67af834b4a00a3e0,64'h635ca4a65037bc0f,
64'ha58e12cb3dfcb235,64'heeae6551b9c25fa1,64'h9660d53ce785a6eb,64'h0000000001000000,
64'h5648e94773770554,64'h38bc97652b54c741,64'he5b26839476fb693,64'hea2b744aec8fa32f,
64'hd173df3571510f4e,64'h4d1d3b1e089317fe,64'h357d520570ee9cff,64'h22a03ac5a37f494a,
64'h2232b9aec8ce93fa,64'hc07b88015eb85552,64'had3c8bdb9c10210f,64'he4421e8e1740a9d6,
64'hcc33aa6490382376,64'h1bedcbd2fbca6eeb,64'h920a40facbc68e3c,64'h3fffbfffc0000000,
64'h8bcee4ee3b19eb5e,64'hfbd8cbd92b76859c,64'hcd625bfe12f1b989,64'h10f31cbf85b4ac62,
64'h86b3220f7b78bc1c,64'h5d309357947e804d,64'hba3da4b625519e39,64'h2e60ca9625a7a426,
64'hc7ea3e234135227d,64'had8d8757deb8ca0b,64'h0cf5f0696940147c,64'h2c6b9494aa06f782,
64'h74b1c25907bf9647,64'hfdd5cca957384bf5,64'hb2cc1aa6fcf0b4de,64'h0000000000200000,
64'h8ac91d286e6ee0ab,64'he71792ebc56a98e9,64'hbcb64d0688edf6d3,64'h3d456e893d91f466,
64'h5a2e7be66e2a21ea,64'h49a3a76381126300,64'h26afaa408e1dd3a0,64'hc4540757f46fe92a,
64'hc44657351919d280,64'hd80f70ff6bd70aab,64'h35a7917b53820422,64'h5c8843d182e8153b,
64'h5986754c5207046f,64'ha37db979bf794dde,64'h9241481ed978d1c8,64'h07fff7fff8000000,
64'h5179dc9d87633d6c,64'h9f7b197aa56ed0b4,64'hf9ac4b7ee25e3732,64'hc21e639730b6958d,
64'h90d664416f6f1784,64'h6ba6126a928fd00a,64'hf747b495e4aa33c8,64'h45cc195284b4f485,
64'h78fd47c40826a450,64'hb5b1b0ea5bd71942,64'h819ebe0cad280290,64'hc58d7291d540def1,
64'h2e96384b00f7f2c9,64'h7fbab994cae7097f,64'h565983549f9e169c,64'h0000000000040000,
64'hb15923a46dcddc16,64'hfce2f25c98ad531e,64'hb796c9a0311dbedb,64'h47a8add0e7b23e8d,
64'hcb45cf7c0dc5443e,64'h093474ec70224c60,64'h04d5f54811c3ba74,64'hd88a80ea3e8dfd26,
64'h1888cae6a3233a50,64'hbb01ee1f4d7ae156,64'hc6b4f22eaa704085,64'hab910879905d02a8,
64'h2b30cea96a40e08e,64'h546fb72ef7ef29bc,64'h12482903db2f1a39,64'h00fffeffff000000,
64'h8a2f3b9330ec67ae,64'h93ef632ed4adda17,64'hdf35896f1c4bc6e7,64'h7843cc728616d2b2,
64'h921acc87adede2f1,64'hcd74c24c9251fa02,64'h1ee8f692bc954679,64'h68b98329f0969e91,
64'h0f1fa8f88104d48a,64'hd6b6361c8b7ae329,64'h1033d7c195a50052,64'hf8b1ae515aa81bdf,
64'he5d2c708801efe5a,64'h2ff75732795ce130,64'h8acb306a13f3c2d4,64'h0000000000008000,
64'h562b24744db9bb83,64'h5f9c5e4b5315aa64,64'hb6f2d9336623b7dc,64'h68f515b9bcf647d2,
64'h5968b9ef41b8a888,64'h01268e9d8e04498c,64'h809abea88238774f,64'h5b11501d07d1bfa5,
64'h0311195cd464674a,64'h57603dc3a9af5c2b,64'h78d69e45754e0811,64'h1572210f320ba055,
64'h456619d4ed481c12,64'h8a8df6e55efde538,64'he249051f9b65e348,64'h001fffdfffe00000,
64'h5145e772261d8cf6,64'h327dec65ba95bb43,64'h3be6b12dc38978dd,64'hcf08798d90c2da57,
64'hf243599015bdbc5f,64'hd9ae9848d24a3f41,64'he3dd1ed17792a8d0,64'hed1730645e12d3d3,
64'hc1e3f51e50209a92,64'hfad6c6c2b16f5c66,64'hc2067af772b4a00b,64'h3f1635ca0b55037c,
64'hdcba58e05003dfcc,64'h05feeae64f2b9c26,64'h9159660cc27e785b,64'h0000000000001000,
64'haac5648de9b73771,64'h8bf38bc8ea62b54d,64'h96de5b25ecc476fc,64'hcd1ea2b6779ec8fb,
64'h0b2d173de8371511,64'h8024d1d331c08932,64'h301357d4f0470eea,64'h6b622a0340fa37f5,
64'hc062232ada8c8cea,64'haaec07b7d535eb86,64'hef1ad3c7cea9c103,64'h62ae44218641740b,
64'hc8acc339dda90383,64'h1151bedcabdfbca7,64'h1c4920a3f36cbc69,64'h0003fffbfffc0000,
64'h4a28bcee04c3b19f,64'ha64fbd8c1752b769,64'h677cd62558712f1c,64'h39e10f3192185b4b,
64'h3e486b31e2b7b78c,64'hfb35d3083a4947e9,64'h1c7ba3da2ef2551a,64'hbda2e60bebc25a7b,
64'hd83c7ea30a041353,64'h5f5ad8d8162deb8d,64'hb840cf5e4e569402,64'h87e2c6b8c16aa070,
64'h9b974b1b8a007bfa,64'h40bfdd5c89e57385,64'hb22b2cc0f84fcf0c,64'h0000000000000200,
64'hf558ac90dd36e6ef,64'h717e7178bd4c56aa,64'h92dbcb643d988ee0,64'hb9a3d4562ef3d920,
64'he165a2e6dd06e2a3,64'hd0049a39a6381127,64'hc6026af9de08e1de,64'h6d6c4540081f46ff,
64'hd80c44649b51919e,64'h555d80f6baa6bd71,64'hbde35a7859d53821,64'hac55c88390c82e82,
64'hb91598669bb52071,64'h222a37db757bf795,64'he38924139e6d978e,64'h00007fff7fff8000,
64'h2945179da0987634,64'hf4c9f7b0a2ea56ee,64'h8cef9ac42b0e25e4,64'ha73c21e592430b6a,
64'h87c90d65bc56f6f2,64'hff66ba60274928fe,64'hc38f747a85de4aa4,64'hb7b45cc0dd784b50,
64'hbb078fd3c140826b,64'h6beb5b1aa2c5bd72,64'hd70819eb09cad281,64'h10fc58d7182d540e,
64'hd372e962b1400f80,64'h6817fbab313cae71,64'h964565979f09f9e2,64'h0000000000000040,
64'h3eab1591fba6dcde,64'hce2fce2e57a98ad6,64'h125b796c87b311dc,64'h17347a8ac5de7b24,
64'hbc2cb45c3ba0dc55,64'h3a00934714c70225,64'h58c04d5efbc11c3c,64'h2dad88a7e103e8e0,
64'h5b01888c536a3234,64'heaabb01df754d7af,64'hf7bc6b4e2b3aa705,64'hd58ab90fb21905d1,
64'hf722b30bf376a40f,64'h644546fb0eaf7ef3,64'h5c71248233cdb2f2,64'h00000fffeffff000,
64'h8528a2f334130ec7,64'h5e993ef5d45d4ade,64'h919df3580561c4bd,64'hd4e7843bf248616e,
64'hd0f921abf78adedf,64'h5fecd74bc4e92520,64'h9871ee8ed0bbc955,64'h16f68b981baf096a,
64'hb760f1f9d828104e,64'hcd7d6b629458b7af,64'hfae1033c81395a51,64'h421f8b1aa305aa82,
64'h1a6e5d2c562801f0,64'hed02ff74862795cf,64'hd2c8acb233e13f3d,64'h0000000000000008,
64'h47d562b1ff74db9c,64'h59c5f9c58af5315b,64'h824b6f2d10f6623c,64'h82e68f50d8bbcf65,
64'h7785968b27741b8b,64'h674012688298e045,64'h8b1809ab5f782388,64'h05b5b114fc207d1c,
64'h8b6031110a6d4647,64'h3d5576039eea9af6,64'h7ef78d69656754e1,64'hfab15721164320bb,
64'h3ee456615e6ed482,64'hac88a8dec1d5efdf,64'hcb8e248f8679b65f,64'h000001fffdfffe00,
64'h30a5145e468261d9,64'h4bd327de7a8ba95c,64'h7233be6aa0ac3898,64'h5a9cf0873e490c2e,
64'h3a1f24355ef15bdc,64'h0bfd9ae9789d24a4,64'h730e3dd17a17792b,64'hc2ded1724375e12e,
64'h56ec1e3efb05020a,64'h39afad6c328b16f6,64'hff5c2066b0272b4b,64'hc843f1629460b551,
64'h034dcba58ac5003e,64'h3da05fee70c4f2ba,64'h7a591595e67c27e8,64'h0000000000000001
};
  //------------------------
  // 512
  //------------------------
  localparam [2*512-1:0][63:0] NTT_GF64_FWD_N512_PHI_L = {
64'hab38bf38115ea62c,64'h705cd1e9bb1779ed,64'h6ce8024cb0531c09,64'h80b6b6221f840fa4,
64'h47aaaec033dd535f,64'hbf562ae382c86418,64'h3591151bb83abdfc,64'h0000003fffbfffc0,
64'h897a64fb4f51752c,64'h4b539e10a7c92186,64'h817fb35caf13a495,64'h585bda2e086ebc26,
64'h4735f5ad465162df,64'hf9087e2b728c16ab,64'hc7b40bfd0e189e58,64'hdfffffff20000001,
64'h956717e6822bd4c6,64'h6e0b9a3cd762ef3e,64'hed9d0048b60a6382,64'h9016d6c3c3f081f5,
64'h28f555d7e67baa6c,64'h17eac55c70590c83,64'h86b222a2f70757c0,64'h00000007fff7fff8,
64'h912f4c9ee9ea2ea6,64'h496a73c1d4f92431,64'h702ff66b35e27493,64'h4b0b7b45810dd785,
64'h28e6beb588ca2c5c,64'hbf210fc4ce5182d6,64'h18f6817fa1c313cb,64'hfbffffff04000001,
64'h52ace2fc90457a99,64'h4dc173475aec5de8,64'hddb3a00856c14c71,64'h7202dad8187e103f,
64'h851eaaba7ccf754e,64'ha2fd58aaee0b2191,64'h10d644545ee0eaf8,64'h00000000fffeffff,
64'h5225e9939d3d45d5,64'he92d4e775a9f2487,64'hae05feccc6bc4e93,64'h69616f685021baf1,
64'h851cd7d63119458c,64'h57e421f859ca305b,64'ha31ed02f5438627a,64'hff7fffff00800001,
64'hea559c5eb208af54,64'h09b82e68eb5d8bbd,64'hfbb674002ad8298f,64'h2e405b5ae30fc208,
64'h50a3d5570f99eeaa,64'hf45fab147dc16433,64'h021ac88a8bdc1d5f,64'h1fffffffffffe000,
64'h6a44bd3213a7a8bb,64'h3d25a9cecb53e491,64'hb5c0bfd8f8d789d3,64'hed2c2dec2a04375f,
64'h90a39afa462328b2,64'haafc843e6b39460c,64'hd463da052a870c50,64'hffefffff00100001,
64'h9d4ab38b564115eb,64'h613705ccbd6bb178,64'h3f76ce7fe55b0532,64'h05c80b6b5c61f841,
64'hca147aaa21f33dd6,64'hbe8bf561efb82c87,64'h20435911317b83ac,64'h03fffffffffffc00,
64'had4897a5a274f518,64'he7a4b538f96a7c93,64'hb6b817fa7f1af13b,64'h3da585bd654086ec,
64'hd214735e88c46517,64'h955f90874d6728c2,64'h1a8c7b40a550e18a,64'hfffdffff00020001,
64'hb3a95670cac822be,64'h0c26e0b997ad762f,64'hc7eed9cf3cab60a7,64'he0b9016c8b8c3f09,
64'h59428f55043e67bb,64'h37d17eac1df70591,64'h84086b21a62f7076,64'h007fffffffffff80,
64'h15a912f4b44e9ea3,64'hbcf496a67f2d4f93,64'hb6d702feafe35e28,64'h87b4b0b72ca810de,
64'h3a428e6bb1188ca3,64'hd2abf21029ace519,64'hc3518f6754aa1c32,64'hffffbfff00004001,
64'h56752acdd9590458,64'h2184dc1712f5aec6,64'h38fddb39c7956c15,64'hfc17202cb17187e2,
64'hab2851ea0087ccf8,64'he6fa2fd4a3bee0b3,64'h50810d63f4c5ee0f,64'h000ffffffffffff0,
64'ha2b5225df689d3d5,64'hb79e92d42fe5a9f3,64'h16dae05fd5fc6bc5,64'h50f69616a595021c,
64'ha74851ccd6231195,64'hfa557e4125359ca4,64'hd86a31ec2a954387,64'hfffff7ff00000801,
64'h0acea559bb2b208b,64'h44309b82a25eb5d9,64'h671fbb66d8f2ad83,64'hdf82e404d62e30fd,
64'h15650a3d4010f99f,64'hbcdf45f9f477dc17,64'h2a1021ac5e98bdc2,64'h0001fffffffffffe,
64'h7456a44b5ed13a7b,64'hb6f3d259e5fcb53f,64'h62db5c0b9abf8d79,64'h8a1ed2c254b2a044,
64'h74e90a393ac46233,64'h9f4aafc7a4a6b395,64'h3b0d463d6552a871,64'hfffffeff00000101,
64'ha159d4aa97656412,64'he886136f744bd6bc,64'hace3f76c3b1e55b1,64'h7bf05c803ac5c620,
64'h22aca14788021f34,64'h379be8bf1e8efb83,64'hc5420434cbd317b9,64'h40003fffc0000000,
64'hae8ad488cbda2750,64'h36de7a4b1cbf96a8,64'hec5b6b809357f1b0,64'h9143da57ca965409,
64'hae9d214687588c47,64'h73e955f89494d673,64'he761a8c6ccaa550f,64'hffffffdf00000021,
64'hd42b3a9492ecac83,64'h9d10c26d6e897ad8,64'hf59c7eeca763cab7,64'h0f7e0b900758b8c4,
64'h84559428710043e7,64'ha6f37d1743d1df71,64'hf8a84085b97a62f8,64'h080007fff8000000,
64'h15d15a91197b44ea,64'h06dbcf496397f2d5,64'h1d8b6d70126afe36,64'hf2287b4a1952ca82,
64'h35d3a428b0eb1189,64'hae7d2abe72929acf,64'h3cec3518b9954aa2,64'hfffffffb00000005,
64'hba856751f25d9591,64'h13a2184dadd12f5b,64'h3eb38fdd74ec7957,64'h81efc17180eb1719,
64'h308ab284ee20087d,64'hf4de6fa2087a3bef,64'h1f150810b72f4c5f,64'h010000ffff000000,
64'hc2ba2b51632f689e,64'h60db79e8cc72fe5b,64'h43b16dadc24d5fc7,64'hde450f68832a5951,
64'he6ba7484361d6232,64'h35cfa557ae52535a,64'hc79d86a25732a955,64'h7fffffff00000001,
64'hf750ace95e4bb2b3,64'ha274430915ba25ec,64'h27d671fb8e9d8f2b,64'hf03df82d501d62e4,
64'h661156503dc40110,64'h3e9bcdf4210f477e,64'h23e2a101f6e5e98c,64'h0020001fffe00000,
64'h58574569ec65ed14,64'hac1b6f3c798e5fcc,64'h28762db59849abf9,64'hfbc8a1ec30654b2b,
64'hdcd74e8fc6c3ac47,64'hc6b9f4aa35ca4a6c,64'h78f3b0d3eae6552b,64'hefffffff00000001,
64'hbeea159c8bc97657,64'h944e8860a2b744be,64'ha4face3ed1d3b1e6,64'h9e07bf052a03ac5d,
64'h0cc22aca07b88022,64'h47d379be4421e8f0,64'h847c541fbedcbd32,64'h00040003fffc0000,
64'h8b0ae8acbd8cbda3,64'h95836de70f31cbfa,64'he50ec5b5d3093580,64'hbf79143ce60ca966,
64'h3b9ae9d1d8d87589,64'h98d73e94c6b9494e,64'haf1e7619dd5ccaa6,64'hfdffffff00000001,
64'h37dd42b371792ecb,64'h5289d10bd456e898,64'h549f59c79a3a763d,64'h73c0f7e04540758c,
64'hc198455880f71005,64'h08fa6f37c8843d1e,64'hd08f8a8337db97a7,64'h000080007fff8000,
64'hb1615d14f7b197b5,64'hd2b06dbc21e63980,64'h1ca1d8b6ba6126b0,64'h57ef22875cc1952d,
64'he7735d395b1b0eb2,64'h531ae7d258d7292a,64'h55e3cec2fbab9955,64'hffbfffff00000001,
64'ha6fba855ce2f25da,64'h0a513a217a8add13,64'h6a93eb3893474ec8,64'h8e781efb88a80eb2,
64'h783308aab01ee201,64'h411f4de6b91087a4,64'h3a11f15046fb72f5,64'h000010000ffff000,
64'h762c2ba23ef632f7,64'h1a560db7843cc730,64'h03943b16d74c24d6,64'h6afde4508b9832a6,
64'hdcee6ba66b6361d7,64'hca635cf98b1ae526,64'h6abc79d7ff75732b,64'hfff7ffff00000001,
64'hd4df7509f9c5e4bc,64'ha14a27438f515ba3,64'h0d527d671268e9d9,64'hd1cf03deb11501d7,
64'hef0661147603dc41,64'h8823e9bc572210f5,64'h67423e29a8df6e5f,64'h0000020001fffe00,
64'h2ec5857427dec65f,64'h034ac1b6f08798e6,64'h407287629ae9849b,64'h4d5fbc89d1730655,
64'h3b9dcd74ad6c6c3b,64'h594c6b9ef1635ca5,64'had578f3a5feeae66,64'hfffeffff00000001,
64'h9a9beea0bf38bc98,64'hb42944e7d1ea2b75,64'he1aa4fac024d1d3c,64'h3a39e07bb622a03b,
64'hfde0cc21aec07b89,64'h71047d372ae4421f,64'h2ce847c5151bedcc,64'h00000040003fffc0,
64'h25d8b0ae64fbd8cc,64'h406958369e10f31d,64'ha80e50ebb35d3094,64'h69abf790da2e60cb,
64'ha773b9adf5ad8d88,64'h6b298d737e2c6b95,64'h55aaf1e70bfdd5cd,64'hffffdfff00000001,
64'h13537dd417e71793,64'h7685289c9a3d456f,64'h9c3549f50049a3a8,64'ha7473c0ed6c45408,
64'hffbc198355d80f72,64'h2e208fa6c55c8844,64'h859d08f822a37dba,64'h000000080007fff8,
64'h84bb16154c9f7b1a,64'h680d2b0673c21e64,64'h9501ca1cf66ba613,64'had357ef17b45cc1a,
64'h14ee7735beb5b1b1,64'h6d6531ae0fc58d73,64'h6ab55e3c817fbaba,64'hfffffbff00000001,
64'ha26a6fb9e2fce2f3,64'h2ed0a5137347a8ae,64'h1386a93ea0093475,64'h14e8e781dad88a81,
64'hdff7832faabb01ef,64'h85c411f458ab9109,64'hd0b3a11e44546fb8,64'h000000010000ffff,
64'hd09762c1e993ef64,64'h8d01a5604e7843cd,64'hb2a03942fecd74c3,64'hd5a6afdd6f68b984,
64'he29dcee5d7d6b637,64'hadaca63521f8b1af,64'hcd56abc6d02ff758,64'hffffff7f00000001,
64'hb44d4df69c5f9c5f,64'h45da14a22e68f516,64'h6270d5277401268f,64'he29d1cef5b5b1151,
64'h3bfef065d557603e,64'hf0b8823dab157222,64'h1a167423c88a8df7,64'h2000000000002000,
64'h9a12ec57bd327ded,64'h71a034aba9cf087a,64'hb6540727bfd9ae99,64'h9ab4d5fb2ded1731,
64'h3c53b9dc9afad6c7,64'h35b594c6843f1636,64'h19aad578da05feeb,64'hffffffef00000001,
64'h3689a9beb38bf38c,64'h48bb429405cd1ea3,64'h2c4e1aa4ce8024d2,64'hfc53a39d0b6b622b,
64'h477fde0c7aaaec08,64'hde171046f562ae45,64'h2342ce84591151bf,64'h0400000000000400,
64'h73425d8a97a64fbe,64'hce340694b539e110,64'hf6ca80e417fb35d4,64'hf3569abe85bda2e7,
64'h278a773b735f5ad9,64'h46b6b2989087e2c7,64'ha3355aae7b40bfde,64'hfffffffd00000001,
64'h86d1353756717e72,64'ha9176851e0b9a3d5,64'hc589c353d9d0049b,64'hbf8a7473016d6c46,
64'h08effbc18f555d81,64'h7bc2e2087eac55c9,64'h246859d06b222a38,64'h0080000000000080,
64'h4e684bb112f4c9f8,64'h19c680d296a73c22,64'h9ed9501c02ff66bb,64'h3e6ad357b0b7b45d,
64'he4f14ee68e6beb5c,64'h28d6d652f210fc59,64'h5466ab558f6817fc,64'hfffffffec0000001,
64'hd0da26a62ace2fcf,64'h7522ed09dc17347b,64'hb8b13869db3a0094,64'h57f14e8e202dad89,
64'he11dff7751eaabb1,64'hef785c402fd58aba,64'h048d0b3a0d644547,64'h0010000000000010,
64'h09cd0976225e993f,64'hc338d01992d4e785,64'hb3db2a02e05fecd8,64'h67cd5a6a9616f68c,
64'h9c9e29dc51cd7d6c,64'he51adac97e421f8c,64'h8a8cd56a31ed0300,64'hfffffffef8000001,
64'h3a1b44d4a559c5fa,64'haea45da09b82e690,64'h9716270cbb674013,64'heafe29d0e405b5b2,
64'hfc23bfee0a3d5577,64'hddef0b8745fab158,64'h2091a16721ac88a9,64'h0002000000000002,
64'h2139a12ea44bd328,64'h78671a02d25a9cf1,64'h167b65405c0bfd9b,64'h8cf9ab4cd2c2ded2,
64'h9393c53b0a39afae,64'h9ca35b58afc843f2,64'h11519aad463da060,64'hfffffffeff000001,
64'hc7436899d4ab38c0,64'h15d48bb413705cd2,64'hb2e2c4e0f76ce803,64'hdd5fc5395c80b6b7,
64'h3f8477fda147aaaf,64'h1bbde170e8bf562b,64'he412342c04359116,64'hc0003fff40000001,
64'h04273425d4897a65,64'hef0ce33f7a4b539f,64'ha2cf6ca76b817fb4,64'hd19f3568da585bdb,
64'h527278a7214735f6,64'hd3946b6a55f9087f,64'h022a3355a8c7b40c,64'hfffffffeffe00001,
64'h18e86d133a956718,64'hc2ba9175c26e0b9b,64'hb65c589b7eed9d01,64'h3babf8a70b9016d7,
64'h27f08eff9428f556,64'ha377bc2d7d17eac6,64'h5c8246854086b223,64'hf80007ff08000001,
64'h6084e6845a912f4d,64'h3de19c67cf496a74,64'h9459ed946d702ff7,64'hba33e6ac7b4b0b7c,
64'h4a4e4f14a428e6bf,64'h3a728d6d2abf2110,64'h8045466a3518f682,64'hfffffffefffc0001,
64'h031d0da26752ace3,64'hb857522e184dc174,64'hf6cb8b128fddb3a1,64'h27757f14c17202db,
64'h44fe11dfb2851eab,64'h546ef7856fa2fd59,64'hab9048d00810d645,64'hff0000ff01000001,
64'h6c109cd02b5225ea,64'h87bc338c79e92d4f,64'h328b3db26dae05ff,64'h97467cd50f696170,
64'h2949c9e274851cd8,64'h074e51ada557e422,64'hd008a8cc86a31ed1,64'hfffffffeffff8001,
64'ha063a1b3acea559d,64'h970aea454309b82f,64'hfed9716171fbb675,64'ha4eeafe1f82e405c,
64'ha89fc23b5650a3d6,64'hea8ddeefcdf45fac,64'h75720919a1021ac9,64'hffe0001f00200001,
64'hcd821399456a44be,64'h30f786716f3d25aa,64'h265167b62db5c0c0,64'h12e8cf9aa1ed2c2e,
64'h0529393c4e90a39b,64'hc0e9ca34f4aafc85,64'hfa011518b0d463db,64'hfffffffefffff001,
64'h740c7436159d4ab4,64'h32e15d4888613706,64'h7fdb2e2bce3f76cf,64'h949dd5fbbf05c80c,
64'h5513f8472aca147b,64'h9d51bbdd79be8bf6,64'heeae41225420435a,64'hfffc000300040001,
64'h59b04272e8ad4898,64'hc61ef0cd6de7a4b6,64'h04ca2cf6c5b6b818,64'h425d19f3143da586,
64'ha0a52726e9d21474,64'h781d39463e955f91,64'hbf4022a2761a8c7c,64'hfffffffefffffe01,
64'h8e818e8642b3a957,64'h465c2ba8d10c26e1,64'h2ffb65c559c7eeda,64'h9293babef7e0b902,
64'haaa27f0845594290,64'h53aa377b6f37d17f,64'hddd5c8238a84086c,64'hffff7fff80008001,
64'h0b36084e5d15a913,64'h58c3de196dbcf497,64'h0099459ed8b6d703,64'h484ba33e2287b4b1,
64'h9414a4e45d3a428f,64'hef03a727e7d2abf3,64'h97e80453cec35190,64'hfffffffeffffffc1,
64'h31d031d0a856752b,64'he8cb85743a2184dd,64'hc5ff6cb7eb38fddc,64'hd25277571efc1721,
64'h15544fe108ab2852,64'h2a7546ef4de6fa30,64'h9bbab903f150810e,64'hffffefff10001001,
64'ha166c1092ba2b523,64'h2b187bc30db79e93,64'ha01328b33b16dae1,64'he9097466e450f697,
64'h3282949c6ba74852,64'hbde074e45cfa557f,64'h12fd008a79d86a32,64'hfffffffefffffff9,
64'ha63a0639750acea6,64'h7d1970ae2744309c,64'h98bfed967d671fbc,64'hfa4a4eea03df82e5,
64'hc2aa89fb6115650b,64'h054ea8dde9bcdf46,64'h537757203e2a1022,64'hfffffdff02000201,
64'hb42cd820857456a5,64'ha5630f77c1b6f3d3,64'hf40265158762db5d,64'h3d212e8cbc8a1ed3,
64'hc6505292cd74e90b,64'h37bc0e9c6b9f4ab0,64'hc25fa0108f3b0d47,64'hffffffff00000000,
64'h54c740c6eea159d5,64'h8fa32e1544e88614,64'h9317fdb24face3f8,64'h7f4949dce07bf05d,
64'hb855513ecc22aca2,64'h40a9d51b7d379be9,64'hca6eeae347c54205,64'hffffffbf00400041,
64'h76859b03b0ae8ad5,64'hb4ac61ee5836de7b,64'h7e804ca250ec5b6c,64'ha7a425d0f79143db,
64'hb8ca0a51b9ae9d22,64'h06f781d38d73e956,64'h384bf401f1e761a9,64'h1fffffffe0000000,
64'h6a98e8187dd42b3b,64'h91f465c2289d10c3,64'h1262ffb649f59c7f,64'h6fe9293b3c0f7e0c,
64'hd70aaa2719845595,64'he8153aa28fa6f37e,64'h794ddd5c08f8a841,64'hfffffff700080009,
64'h6ed0b3601615d15b,64'hb6958c3d2b06dbd0,64'h8fd00993ca1d8b6e,64'hb4f484b97ef2287c,
64'hd71941497735d3a5,64'h40def03a31ae7d2b,64'he7097e7f5e3cec36,64'h03fffffffc000000,
64'had531d026fba8568,64'hb23e8cb7a513a219,64'h224c5ff6a93eb390,64'h8dfd2526e781efc2,
64'h7ae1554483308ab3,64'h5d02a75411f4de70,64'hef29bbaaa11f1509,64'hfffffffe00010002,
64'hadda166b62c2ba2c,64'h16d2b187a560db7a,64'h51fa01323943b16e,64'h969e9096afde4510,
64'h7ae32828cee6ba75,64'ha81bde06a635cfa6,64'h5ce12fcfabc79d87,64'h007fffffff800000,
64'h15aa63a04df750ad,64'hf647d19614a27444,64'h04498bfed527d672,64'hd1bfa4a41cf03df9,
64'haf5c2aa7f0661157,64'h0ba054ea823e9bce,64'hfde537747423e2a2,64'hdfffffff00002001,
64'h95bb42ccec585746,64'hc2da563034ac1b70,64'h4a3f40260728762e,64'h12d3d212d5fbc8a2,
64'h6f5c6504b9dcd74f,64'h55037bc094c6b9f5,64'h2b9c25f9d578f3b1,64'h000ffffffff00000,
64'h62b54c73a9beea16,64'h9ec8fa3242944e89,64'hc089317f1aa4facf,64'hfa37f493a39e07c0,
64'h35eb8554de0cc22b,64'h41740a9d1047d37a,64'hdfbca6edce847c55,64'hfbffffff00000401,
64'h52b768595d8b0ae9,64'h185b4ac60695836e,64'h4947e80480e50ec6,64'hc25a7a419abf7915,
64'h2deb8ca0773b9aea,64'h6aa06f77b298d73f,64'he57384be5aaf1e77,64'h0001fffffffe0000,
64'h4c56a98e3537dd43,64'hf3d91f45685289d2,64'h3811262fc3549f5a,64'h1f46fe927473c0f8,
64'ha6bd70a9fbc19846,64'hc82e8152e208fa70,64'h7bf794dd59d08f8b,64'hff7fffff00000081,
64'hea56ed0a4bb1615e,64'h430b695880d2b06e,64'h4928fd00501ca1d9,64'h784b4f47d357ef23,
64'hc5bd71934ee7735e,64'h2d540deed6531ae8,64'h3cae7097ab55e3cf,64'h00003fffffffc000,
64'ha98ad53126a6fba9,64'hde7b23e7ed0a513b,64'hc70224c5386a93ec,64'h03e8dfd24e8e781f,
64'h54d7ae14ff783309,64'h1905d02a5c411f4e,64'haf7ef29b0b3a11f2,64'hffefffff00000011,
64'h5d4adda109762c2c,64'h48616d2ad01a560e,64'he9251f9f2a03943c,64'haf0969e85a6afde5,
64'h58b7ae3229dcee6c,64'h05aa81bddaca635d,64'h2795ce12d56abc7a,64'h000007fffffff800,
64'hf5315aa544d4df76,64'hbbcf647c5da14a28,64'h98e04498270d527e,64'h207d1bfa29d1cf04,
64'hea9af5c1bfef0662,64'h4320ba050b8823ea,64'hd5efde52a167423f,64'hfffdffff00000003,
64'h8ba95bb3a12ec586,64'h490c2da51a034ac2,64'h9d24a3f365407288,64'h75e12d3cab4d5fbd,
64'h8b16f5c5c53b9dce,64'h60b550375b594c6c,64'hc4f2b9c19aad5790,64'h000000ffffffff00,
64'h5ea62b54689a9bef,64'h1779ec8f8bb42945,64'h531c0892c4e1aa50,64'h840fa37ec53a39e1,
64'hdd535eb777fde0cd,64'hc864173fe171047e,64'h3abdfbca342ce848,64'hbfffbfff40000001,
64'h51752b763425d8b1,64'hc92185b3e3406959,64'h13a4947e6ca80e51,64'h6ebc25a73569abf8,
64'h5162deb878a773ba,64'h8c16aa066b6b298e,64'h189e57383355aaf2,64'h0000001fffffffe0,
64'h2bd4c56a6d13537e,64'h62ef3d9191768529,64'h0a638112589c354a,64'hf081f46ef8a7473d,
64'h7baa6bd68effbc1a,64'h590c82e7bc2e2090,64'h0757bf7946859d09,64'hf7fff7ff08000001,
64'hea2ea56de684bb17,64'hf92430b59c680d2c,64'he274928eed9501cb,64'h0dd784b4e6ad357f,
64'hca2c5bd64f14ee78,64'h5182d5408d6d6532,64'hc313cae6466ab55f,64'h00000003fffffffc,
64'h457a98ad0da26a70,64'hec5de7b1522ed0a6,64'hc14c70218b1386aa,64'h7e103e8d7f14e8e8,
64'hcf754d7a11dff784,64'h0b21905cf785c412,64'he0eaf7ee48d0b3a2,64'hfefffeff01000001,
64'h3d45d4ad9cd09763,64'h9f248616338d01a6,64'hbc4e92513db2a03a,64'h21baf0967cd5a6b0,
64'h19458b7ac9e29dcf,64'hca305aa751adaca7,64'h3862795ca8cd56ac,64'h8000000000000000,
64'h08af5315a1b44d4e,64'h5d8bbcf5ea45da15,64'hd8298e03716270d6,64'h0fc207d1afe29d1d,
64'h99eea9aec23bfef1,64'hc164320adef0b883,64'hdc1d5efd091a1675,64'hffdfffdf00200001,
64'ha7a8ba95139a12ed,64'h53e490c28671a035,64'hd789d24967b65408,64'h04375e12cf9ab4d6,
64'h2328b16f393c53ba,64'h39460b54ca35b595,64'h870c4f2b1519aad6,64'h1000000000000000,
64'h4115ea62743689aa,64'h6bb1779e5d48bb43,64'h5b0531c02e2c4e1b,64'h61f840f9d5fc53a4,
64'hf33dd534f8477fdf,64'hb82c8640bbde1711,64'h7b83abdf412342cf,64'hfffbfffb00040001,
64'h74f517524273425e,64'h6a7c9217f0ce3407,64'h1af13a492cf6ca81,64'h4086ebc219f3569b,
64'hc465162d27278a78,64'h6728c16a3946b6b3,64'h50e189e522a3355b,64'h0200000000000000,
64'hc822bd4b8e86d136,64'had762ef32ba91769,64'hab60a63765c589c4,64'h8c3f081ebabf8a75,
64'h3e67baa67f08effc,64'hf70590c7377bc2e3,64'h2f70757bc824685a,64'hffff7ffe80008001,
64'h4e9ea2ea084e684c,64'h2d4f9242de19c681,64'he35e2748459ed951,64'ha810dd77a33e6ad4,
64'h188ca2c5a4e4f14f,64'hace5182ca728d6d7,64'haa1c313c045466ac,64'h0040000000000000,
64'h590457a931d0da27,64'hf5aec5dd857522ee,64'h956c14c66cb8b139,64'h7187e1037757f14f,
64'h87ccf7544fe11e00,64'hbee0b21846ef785d,64'hc5ee0eaeb9048d0c,64'hffffeffef0001001,
64'h89d3d45cc109cd0a,64'he5a9f2477bc338d1,64'hfc6bc4e828b3db2b,64'h95021bae7467cd5b,
64'h23119458949c9e2a,64'h359ca30574e51adb,64'h95438627008a8cd6,64'h0008000000000000,
64'h2b208af5063a1b45,64'h5eb5d8bb70aea45e,64'hf2ad8297ed971628,64'h2e30fc204eeafe2a,
64'h10f99eea89fc23c0,64'h77dc1642a8ddef0c,64'h98bdc1d5572091a2,64'hfffffdfefe000201,
64'hd13a7a8ad82139a2,64'hfcb53e480f78671b,64'hbf8d789c65167b66,64'hb2a043752e8cf9ac,
64'hc462328a529393c6,64'ha6b394600e9ca35c,64'h52a870c4a011519b,64'h0001000000000000,
64'h6564115e40c74369,64'h4bd6bb172e15d48c,64'h1e55b052fdb2e2c5,64'hc5c61f8349dd5fc6,
64'h021f33dd513f8478,64'h8efb82c7d51bbde2,64'hd317b839eae41235,64'hffffffbeffc00041,
64'hda274f509b042735,64'hbf96a7c861ef0ce4,64'h57f1af134ca2cf6d,64'h9654086e25d19f36,
64'h588c46510a527279,64'h94d6728b81d3946c,64'haa550e17f4022a34,64'h0000200000000000,
64'hecac822ae818e86e,64'h897ad76265c2ba92,64'h63cab609ffb65c59,64'h58b8c3f0293babf9,
64'h0043e67baa27f08f,64'hd1df70583aa377bd,64'h7a62f706dd5c8247,64'hfffffff6fff80009,
64'h7b44e9e9b36084e7,64'h97f2d4f88c3de19d,64'h6afe35e2099459ee,64'h52ca810d84ba33e7,
64'heb1188c9414a4e50,64'h929ace50f03a728e,64'h954aa1c27e804547,64'h0000040000000000,
64'h5d9590451d031d0e,64'hd12f5aeb8cb85753,64'hec7956c05ff6cb8c,64'heb17187d25277580,
64'h20087ccf5544fe12,64'h7a3bee0aa7546ef8,64'h2f4c5ee0bbab9049,64'hfffffffdffff0002,
64'h2f689d3d166c109d,64'h72fe5a9eb187bc34,64'h4d5fc6bc01328b3e,64'h2a5950219097467d,
64'h1d623119282949ca,64'h525359c9de074e52,64'h32a954382fd008a9,64'h0000008000000000,
64'h4bb2b20863a063a2,64'hba25eb5cd1970aeb,64'h9d8f2ad78bfed972,64'h1d62e30fa4a4eeb0,
64'hc4010f992aa89fc3,64'h0f477dc154ea8ddf,64'he5e98bdb3775720a,64'hdffffffeffffe001,
64'h65ed13a742cd8214,64'h8e5fcb535630f787,64'h49abf8d740265168,64'h654b2a03d212e8d0,
64'hc3ac46226505293a,64'hca4a6b387bc0e9cb,64'he6552a8625fa0116,64'h0000001000000000,
64'hc97656404c740c75,64'hb744bd6afa32e15e,64'hd3b1e55a317fdb2f,64'h03ac5c61f4949dd6,
64'hb88021f2855513f9,64'h21e8efb80a9d51bc,64'hdcbd317aa6eeae42,64'hfbfffffefffffc01,
64'h8cbda2746859b043,64'h31cbf96a4ac61ef1,64'h09357f1ae804ca2d,64'h0ca965407a425d1a,
64'hd87588c38ca0a528,64'hb9494d666f781d3a,64'h5ccaa55084bf4023,64'h0000000200000000,
64'h792ecac7a98e818f,64'h56e897ad1f465c2c,64'h3a763cab262ffb66,64'h40758b8bfe9293bb,
64'hf710043d70aaa280,64'h843d1df68153aa38,64'hdb97a62e94ddd5c9,64'hff7ffffeffffff81,
64'hb197b44ded0b3609,64'he6397f2c6958c3df,64'h6126afe2fd009946,64'hc1952ca74f484ba4,
64'h1b0eb118719414a5,64'hd72929ac0def03a8,64'hab9954a97097e805,64'h0000000040000000,
64'h2f25d958d531d032,64'h8add12f523e8cb86,64'h474ec79524c5ff6d,64'ha80eb170dfd25278,
64'h1ee20087ae155450,64'h1087a3bed02a7547,64'hfb72f4c4f29bbaba,64'hffeffffefffffff1,
64'hf632f688dda166c2,64'h3cc72fe56d2b187c,64'h4c24d5fc1fa01329,64'h9832a59469e90975,
64'h6361d622ae328295,64'h1ae5253581bde075,64'h75732a94ce12fd01,64'h0000000008000000,
64'hc5e4bb2a5aa63a07,64'h515ba25e647d1971,64'h68e9d8f24498bfee,64'h1501d62e1bfa4a4f,
64'h03dc4010f5c2aa8a,64'h2210f477ba054ea9,64'hdf6e5e97de537758,64'hfffdfffeffffffff,
64'hdec65ed05bb42cd9,64'h8798e5fc2da56310,64'he9849abea3f40266,64'h730654b22d3d212f,
64'h6c6c3ac3f5c65053,64'h635ca4a65037bc0f,64'heeae6551b9c25fa1,64'h0000000001000000,
64'h38bc97652b54c741,64'hea2b744aec8fa32f,64'h4d1d3b1e089317fe,64'h22a03ac5a37f494a,
64'hc07b88015eb85552,64'he4421e8e1740a9d6,64'h1bedcbd2fbca6eeb,64'h3fffbfffc0000000,
64'hfbd8cbd92b76859c,64'h10f31cbf85b4ac62,64'h5d309357947e804d,64'h2e60ca9625a7a426,
64'had8d8757deb8ca0b,64'h2c6b9494aa06f782,64'hfdd5cca957384bf5,64'h0000000000200000,
64'he71792ebc56a98e9,64'h3d456e893d91f466,64'h49a3a76381126300,64'hc4540757f46fe92a,
64'hd80f70ff6bd70aab,64'h5c8843d182e8153b,64'ha37db979bf794dde,64'h07fff7fff8000000,
64'h9f7b197aa56ed0b4,64'hc21e639730b6958d,64'h6ba6126a928fd00a,64'h45cc195284b4f485,
64'hb5b1b0ea5bd71942,64'hc58d7291d540def1,64'h7fbab994cae7097f,64'h0000000000040000,
64'hfce2f25c98ad531e,64'h47a8add0e7b23e8d,64'h093474ec70224c60,64'hd88a80ea3e8dfd26,
64'hbb01ee1f4d7ae156,64'hab910879905d02a8,64'h546fb72ef7ef29bc,64'h00fffeffff000000,
64'h93ef632ed4adda17,64'h7843cc728616d2b2,64'hcd74c24c9251fa02,64'h68b98329f0969e91,
64'hd6b6361c8b7ae329,64'hf8b1ae515aa81bdf,64'h2ff75732795ce130,64'h0000000000008000,
64'h5f9c5e4b5315aa64,64'h68f515b9bcf647d2,64'h01268e9d8e04498c,64'h5b11501d07d1bfa5,
64'h57603dc3a9af5c2b,64'h1572210f320ba055,64'h8a8df6e55efde538,64'h001fffdfffe00000,
64'h327dec65ba95bb43,64'hcf08798d90c2da57,64'hd9ae9848d24a3f41,64'hed1730645e12d3d3,
64'hfad6c6c2b16f5c66,64'h3f1635ca0b55037c,64'h05feeae64f2b9c26,64'h0000000000001000,
64'h8bf38bc8ea62b54d,64'hcd1ea2b6779ec8fb,64'h8024d1d331c08932,64'h6b622a0340fa37f5,
64'haaec07b7d535eb86,64'h62ae44218641740b,64'h1151bedcabdfbca7,64'h0003fffbfffc0000,
64'ha64fbd8c1752b769,64'h39e10f3192185b4b,64'hfb35d3083a4947e9,64'hbda2e60bebc25a7b,
64'h5f5ad8d8162deb8d,64'h87e2c6b8c16aa070,64'h40bfdd5c89e57385,64'h0000000000000200,
64'h717e7178bd4c56aa,64'hb9a3d4562ef3d920,64'hd0049a39a6381127,64'h6d6c4540081f46ff,
64'h555d80f6baa6bd71,64'hac55c88390c82e82,64'h222a37db757bf795,64'h00007fff7fff8000,
64'hf4c9f7b0a2ea56ee,64'ha73c21e592430b6a,64'hff66ba60274928fe,64'hb7b45cc0dd784b50,
64'h6beb5b1aa2c5bd72,64'h10fc58d7182d540e,64'h6817fbab313cae71,64'h0000000000000040,
64'hce2fce2e57a98ad6,64'h17347a8ac5de7b24,64'h3a00934714c70225,64'h2dad88a7e103e8e0,
64'heaabb01df754d7af,64'hd58ab90fb21905d1,64'h644546fb0eaf7ef3,64'h00000fffeffff000,
64'h5e993ef5d45d4ade,64'hd4e7843bf248616e,64'h5fecd74bc4e92520,64'h16f68b981baf096a,
64'hcd7d6b629458b7af,64'h421f8b1aa305aa82,64'hed02ff74862795cf,64'h0000000000000008,
64'h59c5f9c58af5315b,64'h82e68f50d8bbcf65,64'h674012688298e045,64'h05b5b114fc207d1c,
64'h3d5576039eea9af6,64'hfab15721164320bb,64'hac88a8dec1d5efdf,64'h000001fffdfffe00,
64'h4bd327de7a8ba95c,64'h5a9cf0873e490c2e,64'h0bfd9ae9789d24a4,64'hc2ded1724375e12e,
64'h39afad6c328b16f6,64'hc843f1629460b551,64'h3da05fee70c4f2ba,64'h0000000000000001
};
  //------------------------
  // 256
  //------------------------
  localparam [2*256-1:0][63:0] NTT_GF64_FWD_N256_PHI_L = {
64'h705cd1e9bb1779ed,64'h80b6b6221f840fa4,64'hbf562ae382c86418,64'h0000003fffbfffc0,
64'h4b539e10a7c92186,64'h585bda2e086ebc26,64'hf9087e2b728c16ab,64'hdfffffff20000001,
64'h6e0b9a3cd762ef3e,64'h9016d6c3c3f081f5,64'h17eac55c70590c83,64'h00000007fff7fff8,
64'h496a73c1d4f92431,64'h4b0b7b45810dd785,64'hbf210fc4ce5182d6,64'hfbffffff04000001,
64'h4dc173475aec5de8,64'h7202dad8187e103f,64'ha2fd58aaee0b2191,64'h00000000fffeffff,
64'he92d4e775a9f2487,64'h69616f685021baf1,64'h57e421f859ca305b,64'hff7fffff00800001,
64'h09b82e68eb5d8bbd,64'h2e405b5ae30fc208,64'hf45fab147dc16433,64'h1fffffffffffe000,
64'h3d25a9cecb53e491,64'hed2c2dec2a04375f,64'haafc843e6b39460c,64'hffefffff00100001,
64'h613705ccbd6bb178,64'h05c80b6b5c61f841,64'hbe8bf561efb82c87,64'h03fffffffffffc00,
64'he7a4b538f96a7c93,64'h3da585bd654086ec,64'h955f90874d6728c2,64'hfffdffff00020001,
64'h0c26e0b997ad762f,64'he0b9016c8b8c3f09,64'h37d17eac1df70591,64'h007fffffffffff80,
64'hbcf496a67f2d4f93,64'h87b4b0b72ca810de,64'hd2abf21029ace519,64'hffffbfff00004001,
64'h2184dc1712f5aec6,64'hfc17202cb17187e2,64'he6fa2fd4a3bee0b3,64'h000ffffffffffff0,
64'hb79e92d42fe5a9f3,64'h50f69616a595021c,64'hfa557e4125359ca4,64'hfffff7ff00000801,
64'h44309b82a25eb5d9,64'hdf82e404d62e30fd,64'hbcdf45f9f477dc17,64'h0001fffffffffffe,
64'hb6f3d259e5fcb53f,64'h8a1ed2c254b2a044,64'h9f4aafc7a4a6b395,64'hfffffeff00000101,
64'he886136f744bd6bc,64'h7bf05c803ac5c620,64'h379be8bf1e8efb83,64'h40003fffc0000000,
64'h36de7a4b1cbf96a8,64'h9143da57ca965409,64'h73e955f89494d673,64'hffffffdf00000021,
64'h9d10c26d6e897ad8,64'h0f7e0b900758b8c4,64'ha6f37d1743d1df71,64'h080007fff8000000,
64'h06dbcf496397f2d5,64'hf2287b4a1952ca82,64'hae7d2abe72929acf,64'hfffffffb00000005,
64'h13a2184dadd12f5b,64'h81efc17180eb1719,64'hf4de6fa2087a3bef,64'h010000ffff000000,
64'h60db79e8cc72fe5b,64'hde450f68832a5951,64'h35cfa557ae52535a,64'h7fffffff00000001,
64'ha274430915ba25ec,64'hf03df82d501d62e4,64'h3e9bcdf4210f477e,64'h0020001fffe00000,
64'hac1b6f3c798e5fcc,64'hfbc8a1ec30654b2b,64'hc6b9f4aa35ca4a6c,64'hefffffff00000001,
64'h944e8860a2b744be,64'h9e07bf052a03ac5d,64'h47d379be4421e8f0,64'h00040003fffc0000,
64'h95836de70f31cbfa,64'hbf79143ce60ca966,64'h98d73e94c6b9494e,64'hfdffffff00000001,
64'h5289d10bd456e898,64'h73c0f7e04540758c,64'h08fa6f37c8843d1e,64'h000080007fff8000,
64'hd2b06dbc21e63980,64'h57ef22875cc1952d,64'h531ae7d258d7292a,64'hffbfffff00000001,
64'h0a513a217a8add13,64'h8e781efb88a80eb2,64'h411f4de6b91087a4,64'h000010000ffff000,
64'h1a560db7843cc730,64'h6afde4508b9832a6,64'hca635cf98b1ae526,64'hfff7ffff00000001,
64'ha14a27438f515ba3,64'hd1cf03deb11501d7,64'h8823e9bc572210f5,64'h0000020001fffe00,
64'h034ac1b6f08798e6,64'h4d5fbc89d1730655,64'h594c6b9ef1635ca5,64'hfffeffff00000001,
64'hb42944e7d1ea2b75,64'h3a39e07bb622a03b,64'h71047d372ae4421f,64'h00000040003fffc0,
64'h406958369e10f31d,64'h69abf790da2e60cb,64'h6b298d737e2c6b95,64'hffffdfff00000001,
64'h7685289c9a3d456f,64'ha7473c0ed6c45408,64'h2e208fa6c55c8844,64'h000000080007fff8,
64'h680d2b0673c21e64,64'had357ef17b45cc1a,64'h6d6531ae0fc58d73,64'hfffffbff00000001,
64'h2ed0a5137347a8ae,64'h14e8e781dad88a81,64'h85c411f458ab9109,64'h000000010000ffff,
64'h8d01a5604e7843cd,64'hd5a6afdd6f68b984,64'hadaca63521f8b1af,64'hffffff7f00000001,
64'h45da14a22e68f516,64'he29d1cef5b5b1151,64'hf0b8823dab157222,64'h2000000000002000,
64'h71a034aba9cf087a,64'h9ab4d5fb2ded1731,64'h35b594c6843f1636,64'hffffffef00000001,
64'h48bb429405cd1ea3,64'hfc53a39d0b6b622b,64'hde171046f562ae45,64'h0400000000000400,
64'hce340694b539e110,64'hf3569abe85bda2e7,64'h46b6b2989087e2c7,64'hfffffffd00000001,
64'ha9176851e0b9a3d5,64'hbf8a7473016d6c46,64'h7bc2e2087eac55c9,64'h0080000000000080,
64'h19c680d296a73c22,64'h3e6ad357b0b7b45d,64'h28d6d652f210fc59,64'hfffffffec0000001,
64'h7522ed09dc17347b,64'h57f14e8e202dad89,64'hef785c402fd58aba,64'h0010000000000010,
64'hc338d01992d4e785,64'h67cd5a6a9616f68c,64'he51adac97e421f8c,64'hfffffffef8000001,
64'haea45da09b82e690,64'heafe29d0e405b5b2,64'hddef0b8745fab158,64'h0002000000000002,
64'h78671a02d25a9cf1,64'h8cf9ab4cd2c2ded2,64'h9ca35b58afc843f2,64'hfffffffeff000001,
64'h15d48bb413705cd2,64'hdd5fc5395c80b6b7,64'h1bbde170e8bf562b,64'hc0003fff40000001,
64'hef0ce33f7a4b539f,64'hd19f3568da585bdb,64'hd3946b6a55f9087f,64'hfffffffeffe00001,
64'hc2ba9175c26e0b9b,64'h3babf8a70b9016d7,64'ha377bc2d7d17eac6,64'hf80007ff08000001,
64'h3de19c67cf496a74,64'hba33e6ac7b4b0b7c,64'h3a728d6d2abf2110,64'hfffffffefffc0001,
64'hb857522e184dc174,64'h27757f14c17202db,64'h546ef7856fa2fd59,64'hff0000ff01000001,
64'h87bc338c79e92d4f,64'h97467cd50f696170,64'h074e51ada557e422,64'hfffffffeffff8001,
64'h970aea454309b82f,64'ha4eeafe1f82e405c,64'hea8ddeefcdf45fac,64'hffe0001f00200001,
64'h30f786716f3d25aa,64'h12e8cf9aa1ed2c2e,64'hc0e9ca34f4aafc85,64'hfffffffefffff001,
64'h32e15d4888613706,64'h949dd5fbbf05c80c,64'h9d51bbdd79be8bf6,64'hfffc000300040001,
64'hc61ef0cd6de7a4b6,64'h425d19f3143da586,64'h781d39463e955f91,64'hfffffffefffffe01,
64'h465c2ba8d10c26e1,64'h9293babef7e0b902,64'h53aa377b6f37d17f,64'hffff7fff80008001,
64'h58c3de196dbcf497,64'h484ba33e2287b4b1,64'hef03a727e7d2abf3,64'hfffffffeffffffc1,
64'he8cb85743a2184dd,64'hd25277571efc1721,64'h2a7546ef4de6fa30,64'hffffefff10001001,
64'h2b187bc30db79e93,64'he9097466e450f697,64'hbde074e45cfa557f,64'hfffffffefffffff9,
64'h7d1970ae2744309c,64'hfa4a4eea03df82e5,64'h054ea8dde9bcdf46,64'hfffffdff02000201,
64'ha5630f77c1b6f3d3,64'h3d212e8cbc8a1ed3,64'h37bc0e9c6b9f4ab0,64'hffffffff00000000,
64'h8fa32e1544e88614,64'h7f4949dce07bf05d,64'h40a9d51b7d379be9,64'hffffffbf00400041,
64'hb4ac61ee5836de7b,64'ha7a425d0f79143db,64'h06f781d38d73e956,64'h1fffffffe0000000,
64'h91f465c2289d10c3,64'h6fe9293b3c0f7e0c,64'he8153aa28fa6f37e,64'hfffffff700080009,
64'hb6958c3d2b06dbd0,64'hb4f484b97ef2287c,64'h40def03a31ae7d2b,64'h03fffffffc000000,
64'hb23e8cb7a513a219,64'h8dfd2526e781efc2,64'h5d02a75411f4de70,64'hfffffffe00010002,
64'h16d2b187a560db7a,64'h969e9096afde4510,64'ha81bde06a635cfa6,64'h007fffffff800000,
64'hf647d19614a27444,64'hd1bfa4a41cf03df9,64'h0ba054ea823e9bce,64'hdfffffff00002001,
64'hc2da563034ac1b70,64'h12d3d212d5fbc8a2,64'h55037bc094c6b9f5,64'h000ffffffff00000,
64'h9ec8fa3242944e89,64'hfa37f493a39e07c0,64'h41740a9d1047d37a,64'hfbffffff00000401,
64'h185b4ac60695836e,64'hc25a7a419abf7915,64'h6aa06f77b298d73f,64'h0001fffffffe0000,
64'hf3d91f45685289d2,64'h1f46fe927473c0f8,64'hc82e8152e208fa70,64'hff7fffff00000081,
64'h430b695880d2b06e,64'h784b4f47d357ef23,64'h2d540deed6531ae8,64'h00003fffffffc000,
64'hde7b23e7ed0a513b,64'h03e8dfd24e8e781f,64'h1905d02a5c411f4e,64'hffefffff00000011,
64'h48616d2ad01a560e,64'haf0969e85a6afde5,64'h05aa81bddaca635d,64'h000007fffffff800,
64'hbbcf647c5da14a28,64'h207d1bfa29d1cf04,64'h4320ba050b8823ea,64'hfffdffff00000003,
64'h490c2da51a034ac2,64'h75e12d3cab4d5fbd,64'h60b550375b594c6c,64'h000000ffffffff00,
64'h1779ec8f8bb42945,64'h840fa37ec53a39e1,64'hc864173fe171047e,64'hbfffbfff40000001,
64'hc92185b3e3406959,64'h6ebc25a73569abf8,64'h8c16aa066b6b298e,64'h0000001fffffffe0,
64'h62ef3d9191768529,64'hf081f46ef8a7473d,64'h590c82e7bc2e2090,64'hf7fff7ff08000001,
64'hf92430b59c680d2c,64'h0dd784b4e6ad357f,64'h5182d5408d6d6532,64'h00000003fffffffc,
64'hec5de7b1522ed0a6,64'h7e103e8d7f14e8e8,64'h0b21905cf785c412,64'hfefffeff01000001,
64'h9f248616338d01a6,64'h21baf0967cd5a6b0,64'hca305aa751adaca7,64'h8000000000000000,
64'h5d8bbcf5ea45da15,64'h0fc207d1afe29d1d,64'hc164320adef0b883,64'hffdfffdf00200001,
64'h53e490c28671a035,64'h04375e12cf9ab4d6,64'h39460b54ca35b595,64'h1000000000000000,
64'h6bb1779e5d48bb43,64'h61f840f9d5fc53a4,64'hb82c8640bbde1711,64'hfffbfffb00040001,
64'h6a7c9217f0ce3407,64'h4086ebc219f3569b,64'h6728c16a3946b6b3,64'h0200000000000000,
64'had762ef32ba91769,64'h8c3f081ebabf8a75,64'hf70590c7377bc2e3,64'hffff7ffe80008001,
64'h2d4f9242de19c681,64'ha810dd77a33e6ad4,64'hace5182ca728d6d7,64'h0040000000000000,
64'hf5aec5dd857522ee,64'h7187e1037757f14f,64'hbee0b21846ef785d,64'hffffeffef0001001,
64'he5a9f2477bc338d1,64'h95021bae7467cd5b,64'h359ca30574e51adb,64'h0008000000000000,
64'h5eb5d8bb70aea45e,64'h2e30fc204eeafe2a,64'h77dc1642a8ddef0c,64'hfffffdfefe000201,
64'hfcb53e480f78671b,64'hb2a043752e8cf9ac,64'ha6b394600e9ca35c,64'h0001000000000000,
64'h4bd6bb172e15d48c,64'hc5c61f8349dd5fc6,64'h8efb82c7d51bbde2,64'hffffffbeffc00041,
64'hbf96a7c861ef0ce4,64'h9654086e25d19f36,64'h94d6728b81d3946c,64'h0000200000000000,
64'h897ad76265c2ba92,64'h58b8c3f0293babf9,64'hd1df70583aa377bd,64'hfffffff6fff80009,
64'h97f2d4f88c3de19d,64'h52ca810d84ba33e7,64'h929ace50f03a728e,64'h0000040000000000,
64'hd12f5aeb8cb85753,64'heb17187d25277580,64'h7a3bee0aa7546ef8,64'hfffffffdffff0002,
64'h72fe5a9eb187bc34,64'h2a5950219097467d,64'h525359c9de074e52,64'h0000008000000000,
64'hba25eb5cd1970aeb,64'h1d62e30fa4a4eeb0,64'h0f477dc154ea8ddf,64'hdffffffeffffe001,
64'h8e5fcb535630f787,64'h654b2a03d212e8d0,64'hca4a6b387bc0e9cb,64'h0000001000000000,
64'hb744bd6afa32e15e,64'h03ac5c61f4949dd6,64'h21e8efb80a9d51bc,64'hfbfffffefffffc01,
64'h31cbf96a4ac61ef1,64'h0ca965407a425d1a,64'hb9494d666f781d3a,64'h0000000200000000,
64'h56e897ad1f465c2c,64'h40758b8bfe9293bb,64'h843d1df68153aa38,64'hff7ffffeffffff81,
64'he6397f2c6958c3df,64'hc1952ca74f484ba4,64'hd72929ac0def03a8,64'h0000000040000000,
64'h8add12f523e8cb86,64'ha80eb170dfd25278,64'h1087a3bed02a7547,64'hffeffffefffffff1,
64'h3cc72fe56d2b187c,64'h9832a59469e90975,64'h1ae5253581bde075,64'h0000000008000000,
64'h515ba25e647d1971,64'h1501d62e1bfa4a4f,64'h2210f477ba054ea9,64'hfffdfffeffffffff,
64'h8798e5fc2da56310,64'h730654b22d3d212f,64'h635ca4a65037bc0f,64'h0000000001000000,
64'hea2b744aec8fa32f,64'h22a03ac5a37f494a,64'he4421e8e1740a9d6,64'h3fffbfffc0000000,
64'h10f31cbf85b4ac62,64'h2e60ca9625a7a426,64'h2c6b9494aa06f782,64'h0000000000200000,
64'h3d456e893d91f466,64'hc4540757f46fe92a,64'h5c8843d182e8153b,64'h07fff7fff8000000,
64'hc21e639730b6958d,64'h45cc195284b4f485,64'hc58d7291d540def1,64'h0000000000040000,
64'h47a8add0e7b23e8d,64'hd88a80ea3e8dfd26,64'hab910879905d02a8,64'h00fffeffff000000,
64'h7843cc728616d2b2,64'h68b98329f0969e91,64'hf8b1ae515aa81bdf,64'h0000000000008000,
64'h68f515b9bcf647d2,64'h5b11501d07d1bfa5,64'h1572210f320ba055,64'h001fffdfffe00000,
64'hcf08798d90c2da57,64'hed1730645e12d3d3,64'h3f1635ca0b55037c,64'h0000000000001000,
64'hcd1ea2b6779ec8fb,64'h6b622a0340fa37f5,64'h62ae44218641740b,64'h0003fffbfffc0000,
64'h39e10f3192185b4b,64'hbda2e60bebc25a7b,64'h87e2c6b8c16aa070,64'h0000000000000200,
64'hb9a3d4562ef3d920,64'h6d6c4540081f46ff,64'hac55c88390c82e82,64'h00007fff7fff8000,
64'ha73c21e592430b6a,64'hb7b45cc0dd784b50,64'h10fc58d7182d540e,64'h0000000000000040,
64'h17347a8ac5de7b24,64'h2dad88a7e103e8e0,64'hd58ab90fb21905d1,64'h00000fffeffff000,
64'hd4e7843bf248616e,64'h16f68b981baf096a,64'h421f8b1aa305aa82,64'h0000000000000008,
64'h82e68f50d8bbcf65,64'h05b5b114fc207d1c,64'hfab15721164320bb,64'h000001fffdfffe00,
64'h5a9cf0873e490c2e,64'hc2ded1724375e12e,64'hc843f1629460b551,64'h0000000000000001
};
  //------------------------
  // 128
  //------------------------
  localparam [2*128-1:0][63:0] NTT_GF64_FWD_N128_PHI_L = {
64'h80b6b6221f840fa4,64'h0000003fffbfffc0,64'h585bda2e086ebc26,64'hdfffffff20000001,
64'h9016d6c3c3f081f5,64'h00000007fff7fff8,64'h4b0b7b45810dd785,64'hfbffffff04000001,
64'h7202dad8187e103f,64'h00000000fffeffff,64'h69616f685021baf1,64'hff7fffff00800001,
64'h2e405b5ae30fc208,64'h1fffffffffffe000,64'hed2c2dec2a04375f,64'hffefffff00100001,
64'h05c80b6b5c61f841,64'h03fffffffffffc00,64'h3da585bd654086ec,64'hfffdffff00020001,
64'he0b9016c8b8c3f09,64'h007fffffffffff80,64'h87b4b0b72ca810de,64'hffffbfff00004001,
64'hfc17202cb17187e2,64'h000ffffffffffff0,64'h50f69616a595021c,64'hfffff7ff00000801,
64'hdf82e404d62e30fd,64'h0001fffffffffffe,64'h8a1ed2c254b2a044,64'hfffffeff00000101,
64'h7bf05c803ac5c620,64'h40003fffc0000000,64'h9143da57ca965409,64'hffffffdf00000021,
64'h0f7e0b900758b8c4,64'h080007fff8000000,64'hf2287b4a1952ca82,64'hfffffffb00000005,
64'h81efc17180eb1719,64'h010000ffff000000,64'hde450f68832a5951,64'h7fffffff00000001,
64'hf03df82d501d62e4,64'h0020001fffe00000,64'hfbc8a1ec30654b2b,64'hefffffff00000001,
64'h9e07bf052a03ac5d,64'h00040003fffc0000,64'hbf79143ce60ca966,64'hfdffffff00000001,
64'h73c0f7e04540758c,64'h000080007fff8000,64'h57ef22875cc1952d,64'hffbfffff00000001,
64'h8e781efb88a80eb2,64'h000010000ffff000,64'h6afde4508b9832a6,64'hfff7ffff00000001,
64'hd1cf03deb11501d7,64'h0000020001fffe00,64'h4d5fbc89d1730655,64'hfffeffff00000001,
64'h3a39e07bb622a03b,64'h00000040003fffc0,64'h69abf790da2e60cb,64'hffffdfff00000001,
64'ha7473c0ed6c45408,64'h000000080007fff8,64'had357ef17b45cc1a,64'hfffffbff00000001,
64'h14e8e781dad88a81,64'h000000010000ffff,64'hd5a6afdd6f68b984,64'hffffff7f00000001,
64'he29d1cef5b5b1151,64'h2000000000002000,64'h9ab4d5fb2ded1731,64'hffffffef00000001,
64'hfc53a39d0b6b622b,64'h0400000000000400,64'hf3569abe85bda2e7,64'hfffffffd00000001,
64'hbf8a7473016d6c46,64'h0080000000000080,64'h3e6ad357b0b7b45d,64'hfffffffec0000001,
64'h57f14e8e202dad89,64'h0010000000000010,64'h67cd5a6a9616f68c,64'hfffffffef8000001,
64'heafe29d0e405b5b2,64'h0002000000000002,64'h8cf9ab4cd2c2ded2,64'hfffffffeff000001,
64'hdd5fc5395c80b6b7,64'hc0003fff40000001,64'hd19f3568da585bdb,64'hfffffffeffe00001,
64'h3babf8a70b9016d7,64'hf80007ff08000001,64'hba33e6ac7b4b0b7c,64'hfffffffefffc0001,
64'h27757f14c17202db,64'hff0000ff01000001,64'h97467cd50f696170,64'hfffffffeffff8001,
64'ha4eeafe1f82e405c,64'hffe0001f00200001,64'h12e8cf9aa1ed2c2e,64'hfffffffefffff001,
64'h949dd5fbbf05c80c,64'hfffc000300040001,64'h425d19f3143da586,64'hfffffffefffffe01,
64'h9293babef7e0b902,64'hffff7fff80008001,64'h484ba33e2287b4b1,64'hfffffffeffffffc1,
64'hd25277571efc1721,64'hffffefff10001001,64'he9097466e450f697,64'hfffffffefffffff9,
64'hfa4a4eea03df82e5,64'hfffffdff02000201,64'h3d212e8cbc8a1ed3,64'hffffffff00000000,
64'h7f4949dce07bf05d,64'hffffffbf00400041,64'ha7a425d0f79143db,64'h1fffffffe0000000,
64'h6fe9293b3c0f7e0c,64'hfffffff700080009,64'hb4f484b97ef2287c,64'h03fffffffc000000,
64'h8dfd2526e781efc2,64'hfffffffe00010002,64'h969e9096afde4510,64'h007fffffff800000,
64'hd1bfa4a41cf03df9,64'hdfffffff00002001,64'h12d3d212d5fbc8a2,64'h000ffffffff00000,
64'hfa37f493a39e07c0,64'hfbffffff00000401,64'hc25a7a419abf7915,64'h0001fffffffe0000,
64'h1f46fe927473c0f8,64'hff7fffff00000081,64'h784b4f47d357ef23,64'h00003fffffffc000,
64'h03e8dfd24e8e781f,64'hffefffff00000011,64'haf0969e85a6afde5,64'h000007fffffff800,
64'h207d1bfa29d1cf04,64'hfffdffff00000003,64'h75e12d3cab4d5fbd,64'h000000ffffffff00,
64'h840fa37ec53a39e1,64'hbfffbfff40000001,64'h6ebc25a73569abf8,64'h0000001fffffffe0,
64'hf081f46ef8a7473d,64'hf7fff7ff08000001,64'h0dd784b4e6ad357f,64'h00000003fffffffc,
64'h7e103e8d7f14e8e8,64'hfefffeff01000001,64'h21baf0967cd5a6b0,64'h8000000000000000,
64'h0fc207d1afe29d1d,64'hffdfffdf00200001,64'h04375e12cf9ab4d6,64'h1000000000000000,
64'h61f840f9d5fc53a4,64'hfffbfffb00040001,64'h4086ebc219f3569b,64'h0200000000000000,
64'h8c3f081ebabf8a75,64'hffff7ffe80008001,64'ha810dd77a33e6ad4,64'h0040000000000000,
64'h7187e1037757f14f,64'hffffeffef0001001,64'h95021bae7467cd5b,64'h0008000000000000,
64'h2e30fc204eeafe2a,64'hfffffdfefe000201,64'hb2a043752e8cf9ac,64'h0001000000000000,
64'hc5c61f8349dd5fc6,64'hffffffbeffc00041,64'h9654086e25d19f36,64'h0000200000000000,
64'h58b8c3f0293babf9,64'hfffffff6fff80009,64'h52ca810d84ba33e7,64'h0000040000000000,
64'heb17187d25277580,64'hfffffffdffff0002,64'h2a5950219097467d,64'h0000008000000000,
64'h1d62e30fa4a4eeb0,64'hdffffffeffffe001,64'h654b2a03d212e8d0,64'h0000001000000000,
64'h03ac5c61f4949dd6,64'hfbfffffefffffc01,64'h0ca965407a425d1a,64'h0000000200000000,
64'h40758b8bfe9293bb,64'hff7ffffeffffff81,64'hc1952ca74f484ba4,64'h0000000040000000,
64'ha80eb170dfd25278,64'hffeffffefffffff1,64'h9832a59469e90975,64'h0000000008000000,
64'h1501d62e1bfa4a4f,64'hfffdfffeffffffff,64'h730654b22d3d212f,64'h0000000001000000,
64'h22a03ac5a37f494a,64'h3fffbfffc0000000,64'h2e60ca9625a7a426,64'h0000000000200000,
64'hc4540757f46fe92a,64'h07fff7fff8000000,64'h45cc195284b4f485,64'h0000000000040000,
64'hd88a80ea3e8dfd26,64'h00fffeffff000000,64'h68b98329f0969e91,64'h0000000000008000,
64'h5b11501d07d1bfa5,64'h001fffdfffe00000,64'hed1730645e12d3d3,64'h0000000000001000,
64'h6b622a0340fa37f5,64'h0003fffbfffc0000,64'hbda2e60bebc25a7b,64'h0000000000000200,
64'h6d6c4540081f46ff,64'h00007fff7fff8000,64'hb7b45cc0dd784b50,64'h0000000000000040,
64'h2dad88a7e103e8e0,64'h00000fffeffff000,64'h16f68b981baf096a,64'h0000000000000008,
64'h05b5b114fc207d1c,64'h000001fffdfffe00,64'hc2ded1724375e12e,64'h0000000000000001
};
  //------------------------
  // 64
  //------------------------
  localparam [2*64-1:0][63:0] NTT_GF64_FWD_N64_PHI_L = {
64'h0000003fffbfffc0,64'hdfffffff20000001,64'h00000007fff7fff8,64'hfbffffff04000001,
64'h00000000fffeffff,64'hff7fffff00800001,64'h1fffffffffffe000,64'hffefffff00100001,
64'h03fffffffffffc00,64'hfffdffff00020001,64'h007fffffffffff80,64'hffffbfff00004001,
64'h000ffffffffffff0,64'hfffff7ff00000801,64'h0001fffffffffffe,64'hfffffeff00000101,
64'h40003fffc0000000,64'hffffffdf00000021,64'h080007fff8000000,64'hfffffffb00000005,
64'h010000ffff000000,64'h7fffffff00000001,64'h0020001fffe00000,64'hefffffff00000001,
64'h00040003fffc0000,64'hfdffffff00000001,64'h000080007fff8000,64'hffbfffff00000001,
64'h000010000ffff000,64'hfff7ffff00000001,64'h0000020001fffe00,64'hfffeffff00000001,
64'h00000040003fffc0,64'hffffdfff00000001,64'h000000080007fff8,64'hfffffbff00000001,
64'h000000010000ffff,64'hffffff7f00000001,64'h2000000000002000,64'hffffffef00000001,
64'h0400000000000400,64'hfffffffd00000001,64'h0080000000000080,64'hfffffffec0000001,
64'h0010000000000010,64'hfffffffef8000001,64'h0002000000000002,64'hfffffffeff000001,
64'hc0003fff40000001,64'hfffffffeffe00001,64'hf80007ff08000001,64'hfffffffefffc0001,
64'hff0000ff01000001,64'hfffffffeffff8001,64'hffe0001f00200001,64'hfffffffefffff001,
64'hfffc000300040001,64'hfffffffefffffe01,64'hffff7fff80008001,64'hfffffffeffffffc1,
64'hffffefff10001001,64'hfffffffefffffff9,64'hfffffdff02000201,64'hffffffff00000000,
64'hffffffbf00400041,64'h1fffffffe0000000,64'hfffffff700080009,64'h03fffffffc000000,
64'hfffffffe00010002,64'h007fffffff800000,64'hdfffffff00002001,64'h000ffffffff00000,
64'hfbffffff00000401,64'h0001fffffffe0000,64'hff7fffff00000081,64'h00003fffffffc000,
64'hffefffff00000011,64'h000007fffffff800,64'hfffdffff00000003,64'h000000ffffffff00,
64'hbfffbfff40000001,64'h0000001fffffffe0,64'hf7fff7ff08000001,64'h00000003fffffffc,
64'hfefffeff01000001,64'h8000000000000000,64'hffdfffdf00200001,64'h1000000000000000,
64'hfffbfffb00040001,64'h0200000000000000,64'hffff7ffe80008001,64'h0040000000000000,
64'hffffeffef0001001,64'h0008000000000000,64'hfffffdfefe000201,64'h0001000000000000,
64'hffffffbeffc00041,64'h0000200000000000,64'hfffffff6fff80009,64'h0000040000000000,
64'hfffffffdffff0002,64'h0000008000000000,64'hdffffffeffffe001,64'h0000001000000000,
64'hfbfffffefffffc01,64'h0000000200000000,64'hff7ffffeffffff81,64'h0000000040000000,
64'hffeffffefffffff1,64'h0000000008000000,64'hfffdfffeffffffff,64'h0000000001000000,
64'h3fffbfffc0000000,64'h0000000000200000,64'h07fff7fff8000000,64'h0000000000040000,
64'h00fffeffff000000,64'h0000000000008000,64'h001fffdfffe00000,64'h0000000000001000,
64'h0003fffbfffc0000,64'h0000000000000200,64'h00007fff7fff8000,64'h0000000000000040,
64'h00000fffeffff000,64'h0000000000000008,64'h000001fffdfffe00,64'h0000000000000001
};
  //------------------------
  // 32
  //------------------------
  localparam [2*32-1:0][63:0] NTT_GF64_FWD_N32_PHI_L = {
64'hdfffffff20000001,64'hfbffffff04000001,64'hff7fffff00800001,64'hffefffff00100001,
64'hfffdffff00020001,64'hffffbfff00004001,64'hfffff7ff00000801,64'hfffffeff00000101,
64'hffffffdf00000021,64'hfffffffb00000005,64'h7fffffff00000001,64'hefffffff00000001,
64'hfdffffff00000001,64'hffbfffff00000001,64'hfff7ffff00000001,64'hfffeffff00000001,
64'hffffdfff00000001,64'hfffffbff00000001,64'hffffff7f00000001,64'hffffffef00000001,
64'hfffffffd00000001,64'hfffffffec0000001,64'hfffffffef8000001,64'hfffffffeff000001,
64'hfffffffeffe00001,64'hfffffffefffc0001,64'hfffffffeffff8001,64'hfffffffefffff001,
64'hfffffffefffffe01,64'hfffffffeffffffc1,64'hfffffffefffffff9,64'hffffffff00000000,
64'h1fffffffe0000000,64'h03fffffffc000000,64'h007fffffff800000,64'h000ffffffff00000,
64'h0001fffffffe0000,64'h00003fffffffc000,64'h000007fffffff800,64'h000000ffffffff00,
64'h0000001fffffffe0,64'h00000003fffffffc,64'h8000000000000000,64'h1000000000000000,
64'h0200000000000000,64'h0040000000000000,64'h0008000000000000,64'h0001000000000000,
64'h0000200000000000,64'h0000040000000000,64'h0000008000000000,64'h0000001000000000,
64'h0000000200000000,64'h0000000040000000,64'h0000000008000000,64'h0000000001000000,
64'h0000000000200000,64'h0000000000040000,64'h0000000000008000,64'h0000000000001000,
64'h0000000000000200,64'h0000000000000040,64'h0000000000000008,64'h0000000000000001
};
  //------------------------
  // 16
  //------------------------
  localparam [2*16-1:0][63:0] NTT_GF64_FWD_N16_PHI_L = {
64'hfbffffff04000001,64'hffefffff00100001,64'hffffbfff00004001,64'hfffffeff00000101,
64'hfffffffb00000005,64'hefffffff00000001,64'hffbfffff00000001,64'hfffeffff00000001,
64'hfffffbff00000001,64'hffffffef00000001,64'hfffffffec0000001,64'hfffffffeff000001,
64'hfffffffefffc0001,64'hfffffffefffff001,64'hfffffffeffffffc1,64'hffffffff00000000,
64'h03fffffffc000000,64'h000ffffffff00000,64'h00003fffffffc000,64'h000000ffffffff00,
64'h00000003fffffffc,64'h1000000000000000,64'h0040000000000000,64'h0001000000000000,
64'h0000040000000000,64'h0000001000000000,64'h0000000040000000,64'h0000000001000000,
64'h0000000000040000,64'h0000000000001000,64'h0000000000000040,64'h0000000000000001
};
  //------------------------
  // 8
  //------------------------
  localparam [2*8-1:0][63:0] NTT_GF64_FWD_N8_PHI_L = {
64'hffefffff00100001,64'hfffffeff00000101,64'hefffffff00000001,64'hfffeffff00000001,
64'hffffffef00000001,64'hfffffffeff000001,64'hfffffffefffff001,64'hffffffff00000000,
64'h000ffffffff00000,64'h000000ffffffff00,64'h1000000000000000,64'h0001000000000000,
64'h0000001000000000,64'h0000000001000000,64'h0000000000001000,64'h0000000000000001
};
  //------------------------
  // 4
  //------------------------
  localparam [2*4-1:0][63:0] NTT_GF64_FWD_N4_PHI_L = {
64'hfffffeff00000101,64'hfffeffff00000001,64'hfffffffeff000001,64'hffffffff00000000,
64'h000000ffffffff00,64'h0001000000000000,64'h0000000001000000,64'h0000000000000001
};

  //========================
  // NTT backward
  //========================
  //------------------------
  // 2048
  //------------------------
  localparam [2*2048-1:0][63:0] NTT_GF64_BWD_N2048_PHI_L = {
64'h984ec5194d005735,64'h7a591595e67c27e8,64'he0428bb72ed7342e,64'h3da05fee70c4f2ba,
64'h400a70e5c5f8ce33,64'h034dcba58ac5003e,64'h7b81570ec9c3fb2d,64'hc843f1629460b551,
64'h9b245e0853bb56ce,64'hff5c2066b0272b4b,64'h1aad7e6cc54703a8,64'h39afad6c328b16f6,
64'h30a727ca9e5732bc,64'h56ec1e3efb05020a,64'h027b13b2934dde7c,64'hc2ded1724375e12e,
64'h0ad43edf0692c92c,64'h730e3dd17a17792b,64'ha533c7cb60b307fc,64'h0bfd9ae9789d24a4,
64'h4d459a4a8284e98b,64'h3a1f24355ef15bdc,64'hb79ec87849961fc5,64'h5a9cf0873e490c2e,
64'h675a8e29087cda4a,64'h7233be6aa0ac3898,64'h724187d9d01eef69,64'h4bd327de7a8ba95c,
64'h45c72d9719b3a6b3,64'h30a5145e468261d9,64'h6d782b160a49de19,64'h000001fffdfffe00,
64'hcce3ca95f8f800f1,64'hcb8e248f8679b65f,64'h3e4a26bf7240baba,64'hac88a8dec1d5efdf,
64'h25905f019401e356,64'h3ee456615e6ed482,64'h696bce641c528b1b,64'hfab15721164320bb,
64'h64cfdb5fa5cc9c15,64'h7ef78d69656754e1,64'hb44766c5c7313173,64'h3d5576039eea9af6,
64'h18c77ae98bac4113,64'h8b6031110a6d4647,64'h3691661676209901,64'h05b5b114fc207d1c,
64'h676f89d9da059271,64'h8b1809ab5f782388,64'hce0429153baad8cf,64'h674012688298e045,
64'h7433805d5592e030,64'h7785968b27741b8b,64'h3a3d1ec00d9ec2fe,64'h82e68f50d8bbcf65,
64'ha6d4e45fbdfdcf0c,64'h824b6f2d10f6623c,64'h895a102c6df5fd70,64'h59c5f9c58af5315b,
64'h388e6fcba4e2fa28,64'h47d562b1ff74db9c,64'h66ccad124ac89242,64'h0000000000000008,
64'hc27628ce6802b9a4,64'hd2c8acb233e13f3d,64'h02145dc076b9a169,64'hed02ff74862795cf,
64'h005387302fc67196,64'h1a6e5d2c562801f0,64'hdc0ab8794e1fd965,64'h421f8b1aa305aa82,
64'hd922f0469ddab66c,64'hfae1033c81395a51,64'hd56bf3662a381d40,64'hcd7d6b629458b7af,
64'h85393e55f2b995df,64'hb760f1f9d828104e,64'h13d89d949a6ef3e0,64'h16f68b981baf096a,
64'h56a1f6f834964960,64'h9871ee8ed0bbc955,64'h299e3e6005983fdb,64'h5fecd74bc4e92520,
64'h6a2cd25614274c56,64'hd0f921abf78adedf,64'hbcf643c74cb0fe23,64'hd4e7843bf248616e,
64'h3ad4714b43e6d24d,64'h919df3580561c4bd,64'h920c3ed180f77b45,64'h5e993ef5d45d4ade,
64'h2e396cbacd9d3596,64'h8528a2f334130ec7,64'h6bc158b3524ef0c5,64'h00000fffeffff000,
64'h671e54b5c7c00782,64'h5c71248233cdb2f2,64'hf25135fc9205d5cf,64'h644546fb0eaf7ef3,
64'h2c82f80da00f1aaf,64'hf722b30bf376a40f,64'h4b5e7323e29458d5,64'hd58ab90fb21905d1,
64'h267edb002e64e0a5,64'hf7bc6b4e2b3aa705,64'ha23b363339898b93,64'heaabb01df754d7af,
64'hc63bd74c5d620898,64'h5b01888c536a3234,64'hb48b30b4b104c807,64'h2dad88a7e103e8e0,
64'h3b7c4ed1d02c9385,64'h58c04d5efbc11c3c,64'h702148afdd56c672,64'h3a00934714c70225,
64'ha19c02edac97017d,64'hbc2cb45c3ba0dc55,64'hd1e8f6016cf617ef,64'h17347a8ac5de7b24,
64'h36a72302efee785b,64'h125b796c87b311dc,64'h4ad081676fafeb7c,64'hce2fce2e57a98ad6,
64'hc4737e5e2717d13f,64'h3eab1591fba6dcde,64'h366568955644920d,64'h0000000000000040,
64'h13b146794015cd1a,64'h964565979f09f9e2,64'h10a2ee03b5cd0b48,64'h6817fbab313cae71,
64'h029c39817e338cb0,64'hd372e962b1400f80,64'he055c3d070fecb22,64'h10fc58d7182d540e,
64'hc917823aeed5b35a,64'hd70819eb09cad281,64'hab5f9b3751c0e9fa,64'h6beb5b1aa2c5bd72,
64'h29c9f2b395ccaef4,64'hbb078fd3c140826b,64'h9ec4eca4d3779f00,64'hb7b45cc0dd784b50,
64'hb50fb7c3a4b24afe,64'hc38f747a85de4aa4,64'h4cf1f3012cc1fed7,64'hff66ba60274928fe,
64'h516692b3a13a62ad,64'h87c90d65bc56f6f2,64'he7b21e3f6587f113,64'ha73c21e592430b6a,
64'hd6a38a5b1f369267,64'h8cef9ac42b0e25e4,64'h9061f69007bbda24,64'hf4c9f7b0a2ea56ee,
64'h71cb65d76ce9acaf,64'h2945179da0987634,64'h5e0ac59d92778625,64'h00007fff7fff8000,
64'h38f2a5b13e003c0d,64'he38924139e6d978e,64'h9289afeb902eae71,64'h222a37db757bf795,
64'h6417c06e0078d577,64'hb91598669bb52071,64'h5af3992114a2c6a6,64'hac55c88390c82e82,
64'h33f6d80273270527,64'hbde35a7859d53821,64'h11d9b19ecc4c5c93,64'h555d80f6baa6bd71,
64'h31deba68eb1044ba,64'hd80c44649b51919e,64'ha45985aa88264033,64'h6d6c4540081f46ff,
64'hdbe2768f81649c27,64'hc6026af9de08e1de,64'h810a4581eab6338d,64'hd0049a39a6381127,
64'h0ce0177264b80be3,64'he165a2e6dd06e2a3,64'h8f47b01167b0bf72,64'hb9a3d4562ef3d920,
64'hb53918187f73c2d7,64'h92dbcb643d988ee0,64'h56840b3d7d7f5bde,64'h717e7178bd4c56aa,
64'h239bf2f738be89f2,64'hf558ac90dd36e6ef,64'hb32b44abb2249067,64'h0000000000000200,
64'h9d8a33ca00ae68d0,64'hb22b2cc0f84fcf0c,64'h8517701dae685a40,64'h40bfdd5c89e57385,
64'h14e1cc0bf19c6580,64'h9b974b1b8a007bfa,64'h02ae1e8a87f65909,64'h87e2c6b8c16aa070,
64'h48bc11dd76ad9aca,64'hb840cf5e4e569402,64'h5afcd9bf8e074fcb,64'h5f5ad8d8162deb8d,
64'h4e4f959dae65779f,64'hd83c7ea30a041353,64'hf627652a9bbcf7fc,64'hbda2e60bebc25a7b,
64'ha87dbe22259257eb,64'h1c7ba3da2ef2551a,64'h678f980b660ff6b6,64'hfb35d3083a4947e9,
64'h8b34959f09d31566,64'h3e486b31e2b7b78c,64'h3d90f2022c3f8891,64'h39e10f3192185b4b,
64'hb51c52def9b49332,64'h677cd62558712f1c,64'h830fb4843dded11c,64'ha64fbd8c1752b769,
64'h8e5b2ebe674d6575,64'h4a28bcee04c3b19f,64'hf0562cee93bc3126,64'h0003fffbfffc0000,
64'hc7952d8af001e067,64'h1c4920a3f36cbc69,64'h944d7f6081757384,64'h1151bedcabdfbca7,
64'h20be037303c6abb5,64'hc8acc339dda90383,64'hd79cc90aa516352e,64'h62ae44218641740b,
64'h9fb6c01499382937,64'hef1ad3c7cea9c103,64'h8ecd8cf66262e498,64'haaec07b7d535eb86,
64'h8ef5d348588225cf,64'hc062232ada8c8cea,64'h22cc2d5941320193,64'h6b622a0340fa37f5,
64'hdf13b4820b24e132,64'h301357d4f0470eea,64'h08522c1355b19c64,64'h8024d1d331c08932,
64'h6700bb9325c05f18,64'h0b2d173de8371511,64'h7a3d808f3d85fb8c,64'hcd1ea2b6779ec8fb,
64'ha9c8c0c8fb9e16b3,64'h96de5b25ecc476fc,64'hb42059edebfadeee,64'h8bf38bc8ea62b54d,
64'h1cdf97bac5f44f8f,64'haac5648de9b73771,64'h995a256291248333,64'h0000000000001000,
64'hec519e540573467c,64'h9159660cc27e785b,64'h28bb80f17342d1fc,64'h05feeae64f2b9c26,
64'ha70e605f8ce32c00,64'hdcba58e05003dfcc,64'h1570f4543fb2c848,64'h3f1635ca0b55037c,
64'h45e08eedb56cd64e,64'hc2067af772b4a00b,64'hd7e6cdfe703a7e56,64'hfad6c6c2b16f5c66,
64'h727cacef732bbcf6,64'hc1e3f51e50209a92,64'hb13b295bdde7bfd9,64'hed1730645e12d3d3,
64'h43edf1162c92bf53,64'he3dd1ed17792a8d0,64'h3c7cc05e307fb5ad,64'hd9ae9848d24a3f41,
64'h59a4acfc4e98ab2c,64'hf243599015bdbc5f,64'hec87901261fc4487,64'hcf08798d90c2da57,
64'ha8e296fccda4998b,64'h3be6b12dc38978dd,64'h187da425eef688dc,64'h327dec65ba95bb43,
64'h72d975f73a6b2ba4,64'h5145e772261d8cf6,64'h82b1677b9de18929,64'h001fffdfffe00000,
64'h3ca96c5d800f0332,64'he249051f9b65e348,64'ha26bfb080bab9c1c,64'h8a8df6e55efde538,
64'h05f01b991e355da7,64'h456619d4ed481c12,64'hbce6485b28b1a96a,64'h1572210f320ba055,
64'hfdb600a8c9c149b4,64'h78d69e45754e0811,64'h766c67b7131724bc,64'h57603dc3a9af5c2b,
64'h77ae9a46c4112e74,64'h0311195cd464674a,64'h16616acb09900c97,64'h5b11501d07d1bfa5,
64'hf89da4165927098a,64'h809abea88238774f,64'h4291609aad8ce320,64'h01268e9d8e04498c,
64'h3805dc9c2e02f8bd,64'h5968b9ef41b8a888,64'hd1ec047cec2fdc5d,64'h68f515b9bcf647d2,
64'h4e46064cdcf0b593,64'hb6f2d9336623b7dc,64'ha102cf745fd6f76b,64'h5f9c5e4b5315aa64,
64'he6fcbdd62fa27c78,64'h562b24744db9bb83,64'hcad12b1889241994,64'h0000000000008000,
64'h628cf2a72b9a33d9,64'h8acb306a13f3c2d4,64'h45dc078c9a168fdf,64'h2ff75732795ce130,
64'h3873030167195ffb,64'he5d2c708801efe5a,64'hab87a2a1fd964240,64'hf8b1ae515aa81bdf,
64'h2f04776fab66b26e,64'h1033d7c195a50052,64'hbf366ff981d3f2aa,64'hd6b6361c8b7ae329,
64'h93e5677e995de7ad,64'h0f1fa8f88104d48a,64'h89d94ae3ef3dfec3,64'h68b98329f0969e91,
64'h1f6f88b36495fa96,64'h1ee8f692bc954679,64'he3e602f283fdad67,64'hcd74c24c9251fa02,
64'hcd2567e474c5595e,64'h921acc87adede2f1,64'h643c809a0fe22431,64'h7843cc728616d2b2,
64'h4714b7eb6d24cc53,64'hdf35896f1c4bc6e7,64'hc3ed212f77b446e0,64'h93ef632ed4adda17,
64'h96cbafbcd3595d1d,64'h8a2f3b9330ec67ae,64'h158b3be0ef0c4944,64'h00fffeffff000000,
64'he54b62ed0078198f,64'h12482903db2f1a39,64'h135fd8455d5ce0db,64'h546fb72ef7ef29bc,
64'h2f80dcc8f1aaed38,64'h2b30cea96a40e08e,64'he73242de458d4b4b,64'hab910879905d02a8,
64'hedb0054d4e0a4d99,64'hc6b4f22eaa704085,64'hb3633dbb98b925dd,64'hbb01ee1f4d7ae156,
64'hbd74d2392089739d,64'h1888cae6a3233a50,64'hb30b56584c8064b8,64'hd88a80ea3e8dfd26,
64'hc4ed20b9c9384c49,64'h04d5f54811c3ba74,64'h148b04d76c6718fe,64'h093474ec70224c60,
64'hc02ee4e27017c5e7,64'hcb45cf7c0dc5443e,64'h8f6023ed617ee2e2,64'h47a8add0e7b23e8d,
64'h72303268e785ac96,64'hb796c9a0311dbedb,64'h08167ba7feb7bb53,64'hfce2f25c98ad531e,
64'h37e5eeb87d13e3b9,64'hb15923a46dcddc16,64'h568958ca4920cc9a,64'h0000000000040000,
64'h1467953c5cd19ec5,64'h565983549f9e169c,64'h2ee03c66d0b47ef6,64'h7fbab994cae7097f,
64'hc398180c38caffd7,64'h2e96384b00f7f2c9,64'h5c3d1514ecb211fb,64'hc58d7291d540def1,
64'h7823bb7e5b35936f,64'h819ebe0cad280290,64'hf9b37fd10e9f954b,64'hb5b1b0ea5bd71942,
64'h9f2b3bf8caef3d64,64'h78fd47c40826a450,64'h4eca572379eff614,64'h45cc195284b4f485,
64'hfb7c459b24afd4b0,64'hf747b495e4aa33c8,64'h1f30179b1fed6b31,64'h6ba6126a928fd00a,
64'h692b3f29a62acaea,64'h90d664416f6f1784,64'h21e404d37f112185,64'hc21e639730b6958d,
64'h38a5bf5d69266296,64'hf9ac4b7ee25e3732,64'h1f690981bda236fa,64'h9f7b197aa56ed0b4,
64'hb65d7dea9acae8e4,64'h5179dc9d87633d6c,64'hac59df0778624a20,64'h07fff7fff8000000,
64'h2a5b176f03c0cc71,64'h9241481ed978d1c8,64'h9afec22aeae706d8,64'ha37db979bf794dde,
64'h7c06e6488d5769bf,64'h5986754c5207046f,64'h399216f92c6a5a51,64'h5c8843d182e8153b,
64'h6d802a7170526cc1,64'h35a7917b53820422,64'h9b19ede1c5c92ee3,64'hd80f70ff6bd70aab,
64'heba691ce044b9ce3,64'hc44657351919d280,64'h985ab2c7640325bb,64'hc4540757f46fe92a,
64'h276905d449c26242,64'h26afaa408e1dd3a0,64'ha45826bb6338c7f0,64'h49a3a76381126300,
64'h0177271980be2f32,64'h5a2e7be66e2a21ea,64'h7b011f6f0bf7170c,64'h3d456e893d91f466,
64'h9181934a3c2d64ad,64'hbcb64d0688edf6d3,64'h40b3dd3ff5bdda98,64'he71792ebc56a98e9,
64'hbf2f75c4e89f1dc7,64'h8ac91d286e6ee0ab,64'hb44ac654490664ce,64'h0000000000200000,
64'ha33ca9e2e68cf628,64'hb2cc1aa6fcf0b4de,64'h7701e33785a3f7af,64'hfdd5cca957384bf5,
64'h1cc0c067c657feb2,64'h74b1c25907bf9647,64'he1e8a8a965908fd6,64'h2c6b9494aa06f782,
64'hc11ddbf5d9ac9b75,64'h0cf5f0696940147c,64'hcd9bfe8f74fcaa51,64'had8d8757deb8ca0b,
64'hf959dfca5779eb1c,64'hc7ea3e234135227d,64'h7652b91dcf7fb09e,64'h2e60ca9625a7a426,
64'hdbe22ce0257ea579,64'hba3da4b625519e39,64'hf980bcd8ff6b5988,64'h5d309357947e804d,
64'h4959f9503156574d,64'h86b3220f7b78bc1c,64'h0f20269cf8890c27,64'h10f31cbf85b4ac62,
64'hc52dfaec493314af,64'hcd625bfe12f1b989,64'hfb484c0ded11b7d0,64'hfbd8cbd92b76859c,
64'hb2ebef59d657471b,64'h8bcee4ee3b19eb5e,64'h62cef840c31250fb,64'h3fffbfffc0000000,
64'h52d8bb791e066387,64'h920a40facbc68e3c,64'hd7f6115b573836bc,64'h1bedcbd2fbca6eeb,
64'he03732476abb4df5,64'hcc33aa6490382376,64'hcc90b7ca6352d287,64'he4421e8e1740a9d6,
64'h6c01538e82936605,64'had3c8bdb9c10210f,64'hd8cf6f122e497714,64'hc07b88015eb85552,
64'h5d348e77225ce711,64'h2232b9aec8ce93fa,64'hc2d5963f20192dd4,64'h22a03ac5a37f494a,
64'h3b482ea34e13120f,64'h357d520570ee9cff,64'h22c135e019c63f7b,64'h4d1d3b1e089317fe,
64'h0bb938cc05f17990,64'hd173df3571510f4e,64'hd808fb7b5fb8b85d,64'hea2b744aec8fa32f,
64'h8c0c9a55e16b2564,64'he5b26839476fb693,64'h059eea01adeed4be,64'h38bc97652b54c741,
64'hf97bae2c44f8ee33,64'h5648e94773770554,64'ha25632a74833266b,64'h0000000001000000,
64'h19e54f1c3467b13b,64'h9660d53ce785a6eb,64'hb80f19bf2d1fbd75,64'heeae6551b9c25fa1,
64'he606033e32bff590,64'ha58e12cb3dfcb235,64'h0f4545522c847ea9,64'h635ca4a65037bc0f,
64'h08eedfb4cd64dba2,64'h67af834b4a00a3e0,64'h6cdff481a7e55282,64'h6c6c3ac3f5c65053,
64'hcacefe59bbcf58d9,64'h3f51f12009a913e2,64'hb295c8f17bfd84ed,64'h730654b22d3d212f,
64'hdf1167072bf52bc2,64'hd1ed25b62a8cf1c3,64'hcc05e6cefb5acc39,64'he9849abea3f40266,
64'h4acfca838ab2ba66,64'h3599107fdbc5e0dc,64'h790134e7c4486138,64'h8798e5fc2da56310,
64'h296fd7684998a572,64'h6b12dff6978dcc42,64'hda426076688dbe79,64'hdec65ed05bb42cd9,
64'h975f7ad3b2ba38d3,64'h5e772775d8cf5aec,64'h1677c209189287d5,64'hfffdfffeffffffff,
64'h96c5dbcaf0331c36,64'h905207da5e3471dc,64'hbfb08ae0b9c1b5da,64'hdf6e5e97de537758,
64'h01b9924255da6fa1,64'h619d532a81c11baa,64'h6485be591a969432,64'h2210f477ba054ea9,
64'h600a9c77149b3025,64'h69e45ee1e0810873,64'hc67b7897724bb89a,64'h03dc4010f5c2aa8a,
64'he9a473bb12e73886,64'h1195cd7746749fcf,64'h16acb1ff00c96e9a,64'h1501d62e1bfa4a4f,
64'hda41751b70989077,64'habea902c8774e7f7,64'h1609af01ce31fbd7,64'h68e9d8f24498bfee,
64'h5dc9c6602f8bcc80,64'h8b9ef9b18a887a6a,64'hc047dbe0fdc5c2e2,64'h515ba25e647d1971,
64'h6064d2b30b592b1c,64'h2d9341d13b7db491,64'h2cf7500d6f76a5f0,64'hc5e4bb2a5aa63a07,
64'hcbdd716927c77191,64'hb2474a3d9bb82a9e,64'h12b1953f41993353,64'h0000000008000000,
64'hcf2a78e1a33d89d8,64'hb306a9eb3c2d3754,64'hc078cdfe68fdeba3,64'h75732a94ce12fd01,
64'h303019f895ffac79,64'h2c70965eefe591a3,64'h7a2a2a916423f548,64'h1ae5253581bde075,
64'h4776fda66b26dd10,64'h3d7c1a5d50051efd,64'h66ffa4103f2a940d,64'h6361d622ae328295,
64'h5677f2d3de7ac6c2,64'hfa8f89014d489f0f,64'h94ae4790dfec2763,64'h9832a59469e90975,
64'hf88b383f5fa95e0a,64'h8f692db754678e12,64'h602f367ddad661c2,64'h4c24d5fc1fa01329,
64'h567e541e5595d32e,64'hacc883ffde2f06df,64'hc809a741224309bd,64'h3cc72fe56d2b187c,
64'h4b7ebb434cc52b8f,64'h5896ffb7bc6e620d,64'hd21303b9446df3c2,64'hf632f688dda166c2,
64'hbafbd6a195d1c694,64'hf3b93bb0c67ad75e,64'hb3be1048c4943ea8,64'hffeffffefffffff1,
64'hb62ede5b8198e1ac,64'h82903ed6f1a38edc,64'hfd84570ace0daecb,64'hfb72f4c4f29bbaba,
64'h0dcc9212aed37d08,64'h0cea99570e08dd4d,64'h242df2cbd4b4a18d,64'h1087a3bed02a7547,
64'h0054e3bba4d98125,64'h4f22f71204084395,64'h33dbc4c1925dc4ca,64'h1ee20087ae155450,
64'h4d239ddf9739c429,64'h8cae6bba33a4fe78,64'hb5658ff8064b74d0,64'ha80eb170dfd25278,
64'hd20ba8e184c483b2,64'h5f5481693ba73fb3,64'hb04d780e718fdeb8,64'h474ec79524c5ff6d,
64'hee4e33037c5e63fe,64'h5cf7cd905443d34c,64'h023edf0dee2e170a,64'h8add12f523e8cb86,
64'h0326959b5ac958dd,64'h6c9a0e8adbeda487,64'h67ba806c7bb52f7f,64'h2f25d958d531d032,
64'h5eeb8b4f3e3b8c82,64'h923a51f1ddc154eb,64'h958ca9fa0cc99a98,64'h0000000040000000,
64'h7953c71319ec4eba,64'h98354f5ee169ba9b,64'h03c66ff947ef5d12,64'hab9954a97097e805,
64'h8180cfc5affd63c7,64'h6384b2f87f2c8d17,64'hd151548e211faa3d,64'hd72929ac0def03a8,
64'h3bb7ed355936e87e,64'hebe0d2eb8028f7e7,64'h37fd2084f954a065,64'h1b0eb118719414a5,
64'hb3bf96a0f3d6360e,64'hd47c48116a44f871,64'ha5723c8aff613b14,64'hc1952ca74f484ba4,
64'hc459c201fd4af049,64'h7b496dbea33c708c,64'h0179b3f1d6b30e0d,64'h6126afe2fd009946,
64'hb3f2a0f4acae996e,64'h66442003f17836f3,64'h404d3a0f12184de2,64'he6397f2c6958c3df,
64'h5bf5da1c66295c76,64'hc4b7fdbfe3731066,64'h90981dd0236f9e0a,64'hb197b44ded0b3609,
64'hd7deb511ae8e349b,64'h9dc9dd8d33d6bae9,64'h9df0824b24a1f53b,64'hff7ffffeffffff81,
64'hb176f2e10cc70d5b,64'h1481f6bb8d1c76dc,64'hec22b85d706d7651,64'hdb97a62e94ddd5c9,
64'h6e649095769be840,64'h6754cab87046ea68,64'h216f965fa5a50c67,64'h843d1df68153aa38,
64'h02a71ddd26cc0928,64'h7917b89220421ca6,64'h9ede260d92ee264f,64'hf710043d70aaa280,
64'h691ceefeb9ce2146,64'h65735dd59d27f3bc,64'hab2c7fc5325ba67b,64'h40758b8bfe9293bb,
64'h905d471226241d8a,64'hfaa40b4bdd39fd96,64'h826bc0788c7ef5bb,64'h3a763cab262ffb66,
64'h72719822e2f31fe9,64'he7be6c84a21e9a5e,64'h11f6f86f7170b850,64'h56e897ad1f465c2c,
64'h1934acdad64ac6e8,64'h64d07459df6d2435,64'h3dd40366dda97bf5,64'h792ecac7a98e818f,
64'hf75c5a7bf1dc640e,64'h91d28f92ee0aa754,64'hac654fd4664cd4bc,64'h0000000200000000,
64'hca9e389bcf6275cd,64'hc1aa7afb0b4dd4d4,64'h1e337fca3f7ae890,64'h5ccaa55084bf4023,
64'h0c067e317feb1e34,64'h1c2597c6f96468b5,64'h8a8aa47708fd51e2,64'hb9494d666f781d3a,
64'hddbf69abc9b743ef,64'h5f0697630147bf31,64'hbfe90428caa50327,64'hd87588c38ca0a528,
64'h9dfcb50c9eb1b06b,64'ha3e240915227c382,64'h2b91e45cfb09d89b,64'h0ca965407a425d1a,
64'h22ce1015ea578242,64'hda4b6df819e3845d,64'h0bcd9f8eb5987068,64'h09357f1ae804ca2d,
64'h9f9507aa6574cb6b,64'h322100228bc1b795,64'h0269d07a90c26f0e,64'h31cbf96a4ac61ef1,
64'hdfaed0e5314ae3ae,64'h25bfee051b98832a,64'h84c0ee851b7cf04c,64'h8cbda2746859b043,
64'hbef5a8937471a4d2,64'hee4eec6d9eb5d744,64'hef84125d250fa9d4,64'hfbfffffefffffc01,
64'h8bb7970d66386ad3,64'ha40fb5dc68e3b6e0,64'h6115c2f2836bb281,64'hdcbd317aa6eeae42,
64'h732484aeb4df41fd,64'h3aa655c68237533d,64'h0b7cb2fe2d286337,64'h21e8efb80a9d51bc,
64'h1538eee936604940,64'hc8bdc4940210e52d,64'hf6f1307097713274,64'hb88021f2855513f9,
64'h48e777f8ce710a2d,64'h2b9aeeafe93f9ddd,64'h5963fe2e92dd33d3,64'h03ac5c61f4949dd6,
64'h82ea38953120ec4c,64'hd5205a65e9cfeca9,64'h135e03c863f7add4,64'hd3b1e55a317fdb2f,
64'h938cc11a1798ff45,64'h3df3642c10f4d2e9,64'h8fb7c37b8b85c280,64'hb744bd6afa32e15e,
64'hc9a566d6b2563740,64'h2683a2d1fb6921a5,64'heea01b37ed4bdfa7,64'hc97656404c740c75,
64'hbae2d3e68ee32069,64'h8e947c9b70553a9c,64'h632a7ea83266a5db,64'h0000001000000000,
64'h54f1c4e47b13ae62,64'h0d53d7de5a6ea69a,64'hf19bfe51fbd74480,64'he6552a8625fa0116,
64'h6033f18bff58f1a0,64'he12cbe37cb2345a8,64'h545523bc47ea8f0c,64'hca4a6b387bc0e9cb,
64'hedfb4d644dba1f72,64'hf834bb1a0a3df986,64'hff48214b55281933,64'hc3ac46226505293a,
64'hefe5a868f58d8354,64'h1f12048f913e1c0b,64'h5c8f22e8d84ec4d7,64'h654b2a03d212e8d0,
64'h167080b052bc120f,64'hd25b6fc6cf1c22e2,64'h5e6cfc75acc38340,64'h49abf8d740265168,
64'hfca83d572ba65b54,64'h910801155e0dbca7,64'h134e83d486137870,64'h8e5fcb535630f787,
64'hfd76872f8a571d6a,64'h2dff7029dcc4194f,64'h2607742cdbe7825c,64'h65ed13a742cd8214,
64'hf7ad44a0a38d268b,64'h72776373f5aeba19,64'h7c2092f0287d4e99,64'hdffffffeffffe001,
64'h5dbcb86f31c35694,64'h207daee8471db6fb,64'h08ae17971b5d9405,64'he5e98bdb3775720a,
64'h99242578a6fa0fe5,64'hd532ae3511ba99e7,64'h5be597f1694319b8,64'h0f477dc154ea8ddf,
64'ha9c77749b3024a00,64'h45ee24a610872962,64'hb789838bbb899399,64'hc4010f992aa89fc3,
64'h473bbfc873885166,64'h5cd7758049fceee7,64'hcb1ff17696e99e96,64'h1d62e30fa4a4eeb0,
64'h1751c4ad8907625c,64'ha902d3354e7f6542,64'h9af01e431fbd6ea0,64'h9d8f2ad78bfed972,
64'h9c6608d4bcc7fa24,64'hef9b216187a69747,64'h7dbe1be05c2e13fc,64'hba25eb5cd1970aeb,
64'h4d2b36bb92b1b9fa,64'h341d1690db490d27,64'h7500d9c66a5efd31,64'h4bb2b20863a063a2,
64'hd7169f3977190343,64'h74a3e4df82a9d4dc,64'h1953f54493352ed5,64'h0000008000000000,
64'ha78e2725d89d730e,64'h6a9ebef2d37534d0,64'h8cdff296deba23f9,64'h32a954382fd008a9,
64'h019f8c62fac78cfd,64'h0965f1c5591a2d39,64'ha2a91de43f54785e,64'h525359c9de074e52,
64'h6fda6b296dd0fb89,64'hc1a5d8d751efcc29,64'hfa410a61a940c991,64'h1d623119282949ca,
64'h7f2d434eac6c1a99,64'hf890247c89f0e058,64'he4791748c27626b6,64'h2a5950219097467d,
64'hb384058295e09078,64'h92db7e3c78e1170a,64'hf367e3af661c19fe,64'h4d5fc6bc01328b3e,
64'he541eac05d32da99,64'h884008aef06de534,64'h9a741ea4309bc380,64'h72fe5a9eb187bc34,
64'hebb4398352b8eb49,64'h6ffb814fe620ca77,64'h303ba167df3c12df,64'h2f689d3d166c109d,
64'hbd6a250c1c693451,64'h93bb1ba2ad75d0c5,64'he104978443ea74c5,64'hfffffffdffff0002,
64'hede5c37b8e1ab49e,64'h03ed774338edb7d7,64'h4570bcb8daeca028,64'h2f4c5ee0bbab9049,
64'hc9212bc937d07f24,64'ha99571ae8dd4cf32,64'hdf2cbf8d4a18cdbe,64'h7a3bee0aa7546ef8,
64'h4e3bba5298124ffb,64'h2f71253284394b0e,64'hbc4c1c62dc4c9cc3,64'h20087ccf5544fe12,
64'h39ddfe459c428b2e,64'he6bbac044fe77736,64'h58ff8bbab74cf4aa,64'heb17187d25277580,
64'hba8e256c483b12e0,64'h481699af73fb2a0b,64'hd780f21cfdeb74fc,64'hec7956c05ff6cb8c,
64'he33046a9e63fd11c,64'h7cd90b133d34ba31,64'hedf0df05e1709fdd,64'hd12f5aeb8cb85753,
64'h6959b5de958dcfce,64'ha0e8b487da486937,64'ha806ce3652f7e985,64'h5d9590451d031d0e,
64'hb8b4f9d1b8c81a12,64'ha51f26ff154ea6dd,64'hca9faa2499a976a8,64'h0000040000000000,
64'h3c713933c4eb986b,64'h54f5f7999ba9a67d,64'h66ff94baf5d11fc4,64'h954aa1c27e804547,
64'h0cfc6317d63c67e8,64'h4b2f8e2ac8d169c8,64'h1548ef26faa3c2eb,64'h929ace50f03a728e,
64'h7ed3594e6e87dc45,64'h0d2ec6c08f7e6142,64'hd20853144a064c81,64'heb1188c9414a4e50,
64'hf96a1a786360d4c5,64'hc48123eb4f8702b9,64'h23c8ba4d13b135a9,64'h52ca810d84ba33e7,
64'h9c202c19af0483bb,64'h96dbf1e7c708b84c,64'h9b3f1d8230e0cfe9,64'h6afe35e2099459ee,
64'h2a0f5609e996d4c1,64'h4200457b836f299c,64'hd3a0f52584de1bfc,64'h97f2d4f88c3de19d,
64'h5da1cc2195c75a41,64'h7fdc0a82310653b5,64'h81dd0b3ff9e096f7,64'h7b44e9e9b36084e7,
64'heb512865e349a283,64'h9dd8dd196bae8624,64'h0824bc291f53a621,64'hfffffff6fff80009,
64'h6f2e1be370d5a4e9,64'h1f6bba19c76dbeb8,64'h2b85e5c8d765013e,64'h7a62f706dd5c8247,
64'h49095e4fbe83f91a,64'h4cab8d796ea6798b,64'hf965fc7050c66dea,64'hd1df70583aa377bd,
64'h71ddd296c0927fd6,64'h7b89299521ca586f,64'he260e31be264e613,64'h0043e67baa27f08f,
64'hceeff22de214596f,64'h35dd60297f3bb9a9,64'hc7fc5dd7ba67a54e,64'h58b8c3f0293babf9,
64'hd4712b6741d896fb,64'h40b4cd7d9fd95056,64'hbc0790edef5ba7da,64'h63cab609ffb65c59,
64'h1982355631fe88d9,64'he6c8589ce9a5d185,64'h6f86f8360b84fee1,64'h897ad76265c2ba92,
64'h4acdaef7ac6e7e6d,64'h0745a443d24349b3,64'h403671b797bf4c23,64'hecac822ae818e86e,
64'hc5a7ce92c640d08b,64'h28f937fdaa7536e3,64'h54fd512acd4bb53a,64'h0000200000000000,
64'he389c99f275cc357,64'ha7afbccedd4d33e6,64'h37fca5daae88fe1d,64'haa550e17f4022a34,
64'h67e318beb1e33f40,64'h597c7158468b4e3e,64'haa477937d51e1758,64'h94d6728b81d3946c,
64'hf69aca76743ee225,64'h697636047bf30a10,64'h904298a850326402,64'h588c46510a527279,
64'hcb50d3ca1b06a621,64'h24091f607c3815c2,64'h1e45d2699d89ad47,64'h9654086e25d19f36,
64'he10160d178241dd4,64'hb6df8f423845c25c,64'hd9f8ec1587067f44,64'h57f1af134ca2cf6d,
64'h507ab0504cb6a607,64'h10022bde1b794cde,64'h9d07a93226f0dfda,64'hbf96a7c861ef0ce4,
64'hed0e610eae3ad206,64'hfee0541488329da5,64'h0ee85a03cf04b7b4,64'hda274f509b042735,
64'h5a8943361a4d1411,64'heec6e8cf5d74311c,64'h4125e148fa9d3108,64'hffffffbeffc00041,
64'h7970df1e86ad2745,64'hfb5dd0ce3b6df5c0,64'h5c2f2e47bb2809ef,64'hd317b839eae41235,
64'h484af27ff41fc8ce,64'h655c6bcd7533cc56,64'hcb2fe38986336f49,64'h8efb82c7d51bbde2,
64'h8eee94b90493fead,64'hdc494cac0e52c375,64'h130718e613273091,64'h021f33dd513f8478,
64'h777f917510a2cb72,64'haeeb014cf9ddcd47,64'h3fe2eec3d33d2a6a,64'hc5c61f8349dd5fc6,
64'ha3895b400ec4b7d2,64'h05a66beefeca82ae,64'he03c87747add3ecb,64'h1e55b052fdb2e2c5,
64'hcc11aab18ff446c8,64'h3642c4ee4d2e8c21,64'h7c37c1b35c27f705,64'h4bd6bb172e15d48c,
64'h566d77bf6373f366,64'h3a2d221e921a4d98,64'h01b38dbebdfa6116,64'h6564115e40c74369,
64'h2d3e749c32068452,64'h47c9bfee53a9b717,64'ha7ea89586a5da9ce,64'h0001000000000000,
64'h1c4e4d003ae61ab1,64'h3d7de67bea699f2b,64'hbfe52ed67447f0e7,64'h52a870c4a011519b,
64'h3f18c5f88f19f9fd,64'hcbe38ac4345a71ee,64'h523bc9c3a8f0babb,64'ha6b394600e9ca35c,
64'hb4d653baa1f71121,64'h4bb1b026df98507d,64'h8214c5468193200c,64'hc462328a529393c6,
64'h5a869e56d8353102,64'h2048fb04e1c0ae0f,64'hf22e934cec4d6a38,64'hb2a043752e8cf9ac,
64'h080b0692c120ee99,64'hb6fc7a16c22e12db,64'hcfc760b23833fa1a,64'hbf8d789c65167b66,
64'h83d5828465b53036,64'h80115ef0dbca66f0,64'he83d49953786fecc,64'hfcb53e480f78671b,
64'h6873087c71d69029,64'hf702a0ab4194ed21,64'h7742d01e7825bda0,64'hd13a7a8ad82139a2,
64'hd44a19b2d268a086,64'h76374681eba188d9,64'h092f0a49d4e9883e,64'hfffffdfefe000201,
64'hcb86f8f735693a25,64'hdaee8678db6fadf9,64'he179723fd9404f76,64'h98bdc1d5572091a2,
64'h42579401a0fe466e,64'h2ae35e6ea99e62ad,64'h597f1c52319b7a42,64'h77dc1642a8ddef0c,
64'h7774a5cc249ff564,64'he24a656672961ba2,64'h9838c73099398488,64'h10f99eea89fc23c0,
64'hbbfc8bab85165b8d,64'h77580a6cceee6a33,64'hff17761f99e9534f,64'h2e30fc204eeafe2a,
64'h1c4ada057625be8b,64'h2d335f77f6541570,64'h01e43baad6e9f651,64'hf2ad8297ed971628,
64'h608d55927fa2363a,64'hb216277369746107,64'he1be0d9de13fb825,64'h5eb5d8bb70aea45e,
64'hb36bbdfd1b9f9b2e,64'hd16910f590d26cbf,64'h0d9c6df5efd308b0,64'h2b208af5063a1b45,
64'h69f3a4e29034228f,64'h3e4dff749d4db8b6,64'h3f544ac852ed4e6b,64'h0008000000000000,
64'he2726801d730d588,64'hebef33e0534cf957,64'hff2976b8a23f8733,64'h95438627008a8cd6,
64'hf8c62fc578cfcfe7,64'h5f1c5627a2d38f6a,64'h91de4e1f4785d5d6,64'h359ca30574e51adb,
64'ha6b29dda0fb88903,64'h5d8d8138fcc283e6,64'h10a62a380c99005c,64'h23119458949c9e2a,
64'hd434f2b8c1a9880e,64'h0247d8280e057077,64'h91749a6e626b51b9,64'h95021bae7467cd5b,
64'h40583496090774c8,64'hb7e3d0bb117096d3,64'h7e3b0597c19fd0ca,64'hfc6bc4e828b3db2b,
64'h1eac14272da981ac,64'h008af78ade53377c,64'h41ea4cb0bc37f659,64'he5a9f2477bc338d1,
64'h439843e68eb48145,64'hb81505610ca76901,64'hba1680f6c12decfd,64'h89d3d45cc109cd0a,
64'ha250cd9c9345042a,64'hb1ba34125d0c46c5,64'h4978524ea74c41f0,64'hffffeffef0001001,
64'h5c37c7bfab49d122,64'hd77433ccdb7d6fc2,64'h0bcb9205ca027ba9,64'hc5ee0eaeb9048d0c,
64'h12bca00f07f2336e,64'h571af3764cf31567,64'hcbf8e2938cdbd20e,64'hbee0b21846ef785d,
64'hbba52e6424ffab1d,64'h12532b3a94b0dd09,64'hc1c63988c9cc243c,64'h87ccf7544fe11e00,
64'hdfe45d6128b2dc63,64'hbac0536977735195,64'hf8bbb103cf4a9a71,64'h7187e1037757f14f,
64'he256d02bb12df458,64'h699afbc0b2a0ab7f,64'h0f21dd56b74fb288,64'h956c14c66cb8b139,
64'h046aac96fd11b1cd,64'h90b13ba04ba30833,64'h0df06cf609fdc121,64'hf5aec5dd857522ee,
64'h9b5defeddcfcd96b,64'h8b4887b2869365f2,64'h6ce36faf7e984580,64'h590457a931d0da27,
64'h4f9d271781a11475,64'hf26ffba5ea6dc5af,64'hfaa25643976a7357,64'h0040000000000000,
64'h13934015b986ac39,64'h5f799f099a67cab1,64'hf94bb5cc11fc3991,64'haa1c313c045466ac,
64'hc6317e32c67e7f31,64'hf8e2b13f169c7b4e,64'h8ef270fe3c2eaeac,64'hace5182ca728d6d7,
64'h3594eed57dc44813,64'hec6c09c9e6141f2e,64'h853151c064c802e0,64'h188ca2c5a4e4f14f,
64'ha1a795cc0d4c406a,64'h123ec140702b83b8,64'h8ba4d377135a8dc4,64'ha810dd77a33e6ad4,
64'h02c1a4b2483ba63e,64'hbf1e85dd8b84b693,64'hf1d82cc10cfe864d,64'he35e2748459ed951,
64'hf560a1396d4c0d60,64'h0457bc56f299bbe0,64'h0f526587e1bfb2c6,64'h2d4f9242de19c681,
64'h1cc21f3675a40a26,64'hc0a82b0d653b4803,64'hd0b407bb096f67e3,64'h4e9ea2ea084e684c,
64'h12866ce99a28214b,64'h8dd1a097e8623623,64'h4bc292773a620f7e,64'hffff7ffe80008001,
64'he1be3dff5a4e890e,64'hbba19e6cdbeb7e0a,64'h5e5c902e5013dd48,64'h2f70757bc824685a,
64'h95e500783f919b70,64'hb8d79bb46798ab36,64'h5fc714a266de906a,64'hf70590c7377bc2e3,
64'hdd29732627fd58e3,64'h929959d4a586e848,64'h0e31cc4c4e6121da,64'h3e67baa67f08effc,
64'hff22eb0f4596e312,64'hd6029b50bb9a8ca3,64'hc5dd88257a54d381,64'h8c3f081ebabf8a75,
64'h12b68164896fa2b9,64'h4cd7de0895055bf5,64'h790eeab5ba7d9440,64'hab60a63765c589c4,
64'h235564b7e88d8e68,64'h8589dd065d184194,64'h6f8367b04fee0908,64'had762ef32ba91769,
64'hdaef7f72e7e6cb54,64'h5a443d98349b2f8c,64'h671b7d7ef4c22bfd,64'hc822bd4b8e86d136,
64'h7ce938be0d08a3a6,64'h937fdd36536e2d71,64'hd512b223bb539ab1,64'h0200000000000000,
64'h9c9a00adcc3561c8,64'hfbccf84ed33e5586,64'hca5dae678fe1cc81,64'h50e189e522a3355b,
64'h318bf19c33f3f982,64'hc71589ffb4e3da69,64'h779387f5e175755c,64'h6728c16a3946b6b3,
64'haca776acee224097,64'h63604e5630a0f969,64'h298a8e07264016fc,64'hc465162d27278a78,
64'h0d3cae656a62034b,64'h91f60a03815c1dc0,64'h5d269bbc9ad46e1c,64'h4086ebc219f3569b,
64'h160d259241dd31f0,64'hf8f42ef15c25b493,64'h8ec1660f67f43261,64'h1af13a492cf6ca81,
64'hab0509d26a606af9,64'h22bde2b794cddf00,64'h7a932c3f0dfd9630,64'h6a7c9217f0ce3407,
64'he610f9b3ad205130,64'h0541587129da4012,64'h85a03dde4b7b3f12,64'h74f517524273425e,
64'h9433674cd1410a58,64'h6e8d04c34311b114,64'h5e1493bbd3107bee,64'hfffbfffb00040001,
64'h0df1f001d2744869,64'hdd0cf36bdf5bf04b,64'hf2e48174809eea3e,64'h7b83abdf412342cf,
64'haf2803c5fc8cdb7c,64'hc6bcdda83cc559ab,64'hfe38a51536f4834e,64'hb82c8640bbde1711,
64'he94b99373feac712,64'h94cacea92c37423c,64'h718e626273090ed0,64'hf33dd534f8477fdf,
64'hf91758812cb71889,64'hb014da8bdcd46512,64'h2eec4131d2a69c02,64'h61f840f9d5fc53a4,
64'h95b40b244b7d15c8,64'h66bef046a82adfa6,64'hc87755b0d3eca1fd,64'h5b0531c02e2c4e1b,
64'h1aab25c0446c733f,64'h2c4ee836e8c20c9c,64'h7c1b3d857f70483d,64'h6bb1779e5d48bb43,
64'hd77bfb9d3f365a9a,64'hd221ecc3a4d97c5e,64'h38dbebfaa6115fe5,64'h4115ea62743689aa,
64'he749c5f368451d2d,64'h9bfee9b69b716b84,64'ha8959123da9cd582,64'h1000000000000000,
64'he4d0057261ab0e3c,64'hde67c27d99f2ac29,64'h52ed73427f0e6402,64'h870c4f2b1519aad6,
64'h8c5f8ce29f9fcc0f,64'h38ac5003a71ed342,64'hbc9c3fb20babaadd,64'h39460b54ca35b595,
64'h653bb56c711204b3,64'h1b0272b48507cb45,64'h4c54703a3200b7df,64'h2328b16f393c53ba,
64'h69e5732b53101a58,64'h8fb050200ae0edfc,64'he934dde6d6a370de,64'h04375e12cf9ab4d6,
64'hb0692c920ee98f80,64'hc7a17791e12da491,64'h760b307f3fa19304,64'hd789d24967b65408,
64'h58284e98530357c3,64'h15ef15bda66ef7ff,64'hd49961fb6fecb17d,64'h53e490c28671a035,
64'h3087cda469028979,64'h2a0ac3894ed20090,64'h2d01eef65bd9f88c,64'ha7a8ba95139a12ed,
64'ha19b3a6a8a0852bc,64'h7468261d188d889d,64'hf0a49de09883df6e,64'hffdfffdf00200001,
64'h6f8f800e93a24348,64'he8679b64fadf8252,64'h97240bab04f751e9,64'hdc1d5efd091a1675,
64'h79401e34e466dbdb,64'h35e6ed47e62acd52,64'hf1c528b0b7a41a69,64'hc164320adef0b883,
64'h4a5cc9c0ff563889,64'ha656754d61ba11dc,64'h8c7313169848767d,64'h99eea9aec23bfef1,
64'hc8bac41065b8c441,64'h80a6d463e6a3288b,64'h7762098f9534e00f,64'h0fc207d1afe29d1d,
64'hada059265be8ae3c,64'h35f782384156fd2d,64'h43baad8c9f650fe2,64'hd8298e03716270d6,
64'hd5592e02236399f8,64'h627741b8461064df,64'he0d9ec2efb8241e5,64'h5d8bbcf5ea45da15,
64'hbbdfdceff9b2d4ca,64'h910f662326cbe2ea,64'hc6df5fd6308aff27,64'h08af5315a1b44d4e,
64'h3a4e2fa24228e961,64'hdff74db8db8b5c1c,64'h44ac8923d4e6ac0b,64'h8000000000000000,
64'h26802b9a0d5871d9,64'hf33e13f2cf956142,64'h976b9a15f873200e,64'h3862795ca8cd56ac,
64'h62fc6718fcfe6074,64'hc562801e38f69a0f,64'he4e1fd955d5d56e3,64'hca305aa751adaca7,
64'h29ddab6688902595,64'hd81395a4283e5a28,64'h62a381d39005bef6,64'h19458b7ac9e29dcf,
64'h4f2b995d9880d2bd,64'h7d82810457076fdc,64'h49a6ef3db51b86e9,64'h21baf0967cd5a6b0,
64'h83496495774c7bfb,64'h3d0bbc95096d2482,64'hb05983fcfd0c981d,64'hbc4e92513db2a03a,
64'hc14274c4981abe16,64'haf78aded3377bff8,64'ha4cb0fe17f658be2,64'h9f248616338d01a6,
64'h843e6d2448144bc7,64'h50561c4b7690047f,64'h680f77b3decfc45f,64'h3d45d4ad9cd09763,
64'h0cd9d359504295db,64'ha34130ebc46c44e5,64'h8524ef0bc41efb69,64'hfefffeff01000001,
64'h7c7c00779d121a3d,64'h433cdb2ed6fc1289,64'hb9205d5c27ba8f44,64'he0eaf7ee48d0b3a2,
64'hca00f1aa2336ded5,64'haf376a4031566a8f,64'h8e29458cbd20d341,64'h0b21905cf785c412,
64'h52e64e09fab1c446,64'h32b3aa700dd08edb,64'h639898b8c243b3e4,64'hcf754d7a11dff784,
64'h45d620892dc62202,64'h0536a32335194454,64'hbb104c7fa9a70075,64'h7e103e8d7f14e8e8,
64'h6d02c937df4571db,64'hafbc11c30ab7e967,64'h1dd56c66fb287f0e,64'hc14c70218b1386aa,
64'haac970171b1ccfba,64'h13ba0dc5308326f5,64'h06cf617edc120f21,64'hec5de7b1522ed0a6,
64'hdefee784cd96a64b,64'h887b311d365f174c,64'h36fafeb78457f932,64'h457a98ad0da26a70,
64'hd2717d1311474b07,64'hffba6dccdc5ae0da,64'h25644920a7356056,64'h00000003fffffffc,
64'h34015cd16ac38ec7,64'h99f09f9d7cab0a09,64'hbb5cd0b3c399006c,64'hc313cae6466ab55f,
64'h17e338cae7f3039d,64'h2b1400f7c7b4d072,64'h270fecb1eaeab711,64'h5182d5408d6d6532,
64'h4eed5b3544812ca7,64'hc09cad2741f2d13a,64'h151c0e9f802df7ad,64'hca2c5bd64f14ee78,
64'h795ccaeec40695e6,64'hec140825b83b7edd,64'h4d3779efa8dc3746,64'h0dd784b4e6ad357f,
64'h1a4b24afba63dfd4,64'he85de4a94b69240f,64'h82cc1fece864c0e3,64'he274928eed9501cb,
64'h0a13a62ac0d5f0aa,64'h7bc56f6e9bbdffbb,64'h26587f10fb2c5f0b,64'hf92430b59c680d2c,
64'h21f3692640a25e34,64'h82b0e25db48023f6,64'h407bbda1f67e22f5,64'hea2ea56de684bb17,
64'h66ce9aca8214aed8,64'h1a09876323622723,64'h2927786220f7db44,64'hf7fff7ff08000001,
64'he3e003bfe890d1e5,64'h19e6d978b7e09446,64'hc902eae63dd47a1b,64'h0757bf7946859d09,
64'h50078d5719b6f6a2,64'h79bb52068ab35473,64'h714a2c69e9069a04,64'h590c82e7bc2e2090,
64'h97327051d58e222e,64'h959d53816e8476d7,64'h1cc4c5c9121d9f1d,64'h7baa6bd68effbc1a,
64'h2eb1044b6e31100e,64'h29b51919a8ca22a0,64'hd88264024d3803a3,64'hf081f46ef8a7473d,
64'h681649c1fa2b8ed5,64'h7de08e1d55bf4b33,64'heeab6337d943f870,64'h0a638112589c354a,
64'h564b80bdd8e67dcb,64'h9dd06e29841937a8,64'h367b0bf6e0907908,64'h62ef3d9191768529,
64'hf7f73c2c6cb53252,64'h43d988edb2f8ba5c,64'hb7d7f5bd22bfc98f,64'h2bd4c56a6d13537e,
64'h938be89e8a3a5832,64'hfdd36e6de2d706c9,64'h2b22490639ab02af,64'h0000001fffffffe0,
64'ha00ae68c561c7637,64'hcf84fcefe5585044,64'hdae685a31cc8035b,64'h189e57383355aaf2,
64'hbf19c6573f981ce8,64'h58a007bf3da6838f,64'h387f65905755b887,64'h8c16aa066b6b298e,
64'h776ad9ac24096536,64'h04e569400f9689ca,64'ha8e074fc016fbd68,64'h5162deb878a773ba,
64'hcae657792034af2d,64'h60a04134c1dbf6e1,64'h69bbcf7f46e1ba2e,64'h6ebc25a73569abf8,
64'hd259257dd31efea0,64'h42ef25515b492071,64'h1660ff6b43260714,64'h13a4947e6ca80e51,
64'h509d315606af8550,64'hde2b7b77ddeffdd5,64'h32c3f888d962f857,64'hc92185b3e3406959,
64'h0f9b49330512f19f,64'h158712f1a4011fac,64'h03dded11b3f117a6,64'h51752b763425d8b1,
64'h3674d65710a576bd,64'hd04c3b191b113918,64'h493bc31207beda1f,64'hbfffbfff40000001,
64'h1f001e0644868f21,64'hcf36cbc5bf04a230,64'h48175737eea3d0d2,64'h3abdfbca342ce848,
64'h803c6abacdb7b50e,64'hcdda9037559aa395,64'h8a5163524834d01d,64'hc864173fe171047e,
64'hb9938292ac71116c,64'hacea9c0f7423b6b4,64'he6262e4890ecf8e8,64'hdd535eb777fde0cd,
64'h7588225c7188806f,64'h4da8c8ce465114ff,64'hc413201869c01d12,64'h840fa37ec53a39e1,
64'h40b24e12d15c76a5,64'hef0470edadfa5995,64'h755b19c5ca1fc379,64'h531c0892c4e1aa50,
64'hb25c05f0c733ee56,64'hee83715020c9bd3c,64'hb3d85fb80483c83f,64'h1779ec8f8bb42945,
64'hbfb9e16a65a99289,64'h1ecc476f97c5d2de,64'hbebfadee15fe4c73,64'h5ea62b54689a9bef,
64'h9c5f44f851d2c18c,64'hee9b737616b83641,64'h59124832cd581577,64'h000000ffffffff00,
64'h00573467b0e3b1b3,64'h7c27e7852ac2821a,64'hd7342d1ee6401ad2,64'hc4f2b9c19aad5790,
64'hf8ce32befcc0e73b,64'hc5003dfbed341c76,64'hc3fb2c83baadc437,64'h60b550375b594c6c,
64'hbb56cd64204b29ad,64'h272b4a007cb44e50,64'h4703a7e50b7deb3b,64'h8b16f5c5c53b9dce,
64'h5732bbcf01a57962,64'h050209a90edfb705,64'h4dde7bfd370dd16d,64'h75e12d3cab4d5fbd,
64'h92c92bf498f7f4fa,64'h17792a8cda490386,64'hb307fb5a193038a0,64'h9d24a3f365407288,
64'h84e98ab2357c2a7e,64'hf15bdbc4ef7feea2,64'h961fc447cb17c2b7,64'h490c2da51a034ac2,
64'h7cda499828978cf8,64'hac38978d2008fd60,64'h1eef688d9f88bd30,64'h8ba95bb3a12ec586,
64'hb3a6b2b9852bb5e7,64'h8261d8ced889c8ba,64'h49de18923df6d0f6,64'hfffdffff00000003,
64'hf800f03224347908,64'h79b65e33f825117a,64'h40bab9c1751e868e,64'hd5efde52a167423f,
64'h01e355da6dbda86c,64'h6ed481c0acd51ca2,64'h528b1a9641a680e4,64'h4320ba050b8823ea,
64'hcc9c149a63888b5b,64'h6754e080a11db59b,64'h3131724b8767c739,64'hea9af5c1bfef0662,
64'hac4112e68c440375,64'h6d4646743288a7f6,64'h209900c94e00e88a,64'h207d1bfa29d1cf04,
64'h059270988ae3b526,64'h782387746fd2cca1,64'haad8ce3150fe1bc5,64'h98e04498270d527e,
64'h92e02f8b399f72ab,64'h741b8a88064de9d9,64'h9ec2fdc5241e41f3,64'hbbcf647c5da14a28,
64'hfdcf0b582d4c9443,64'hf6623b7cbe2e96f0,64'hf5fd6f75aff26393,64'hf5315aa544d4df76,
64'he2fa27c68e960c5c,64'h74db9bb7b5c1b201,64'hc89241986ac0abb6,64'h000007fffffff800,
64'h02b9a33d871d8d98,64'he13f3c2c561410cd,64'hb9a168fd3200d68a,64'h2795ce12d56abc7a,
64'hc67195fee60739d1,64'h2801efe569a0e3aa,64'h1fd96423d56e21b2,64'h05aa81bddaca635d,
64'hdab66b2602594d63,64'h395a5004e5a2727f,64'h381d3f2a5bef59d6,64'h58b7ae3229dcee6c,
64'hb995de7a0d2bcb0e,64'h28104d4876fdb828,64'h6ef3dfebb86e8b66,64'haf0969e85a6afde5,
64'h96495fa8c7bfa7cc,64'hbbc95466d2481c30,64'h983fdad5c981c4fb,64'he9251f9f2a03943c,
64'h274c5595abe153ec,64'h8adede2e7bff7509,64'hb0fe224258be15b4,64'h48616d2ad01a560e,
64'he6d24cc444bc67bd,64'h61c4bc6e0047eafb,64'hf77b446cfc45e980,64'h5d4adda109762c2c,
64'h9d3595d1295daf33,64'h130ec67ac44e45cc,64'h4ef0c493efb687ae,64'hffefffff00000011,
64'hc007819821a3c839,64'hcdb2f1a2c1288bcd,64'h05d5ce0da8f4346e,64'haf7ef29b0b3a11f2,
64'h0f1aaed36ded4360,64'h76a40e0866a8e50d,64'h9458d4b40d34071e,64'h1905d02a5c411f4e,
64'h64e0a4d91c445ad2,64'h3aa7040808edacd5,64'h898b925d3b3e39c7,64'h54d7ae14ff783309,
64'h6208973962201ba3,64'h6a3233a494453fad,64'h04c8064b7007444f,64'h03e8dfd24e8e781f,
64'h2c9384c4571da930,64'hc11c3ba67e966505,64'h56c6718f87f0de23,64'hc70224c5386a93ec,
64'h97017c5dccfb9554,64'ha0dc5443326f4ec5,64'hf617ee2d20f20f94,64'hde7b23e7ed0a513b,
64'hee785ac86a64a211,64'hb311dbecf174b779,64'hafeb7bb47f931c91,64'ha98ad53126a6fba9,
64'h17d13e3b74b062d9,64'ha6dcddc0ae0d9005,64'h44920cc956055daa,64'h00003fffffffc000,
64'h15cd19ec38ec6cc0,64'h09f9e169b0a08661,64'hcd0b47ee9006b44b,64'h3cae7097ab55e3cf,
64'h338caffd3039ce82,64'h400f7f2c4d071d4f,64'hfecb211eab710d90,64'h2d540deed6531ae8,
64'hd5b3593612ca6b12,64'hcad280282d1393f7,64'hc0e9f953df7aceaf,64'hc5bd71934ee7735e,
64'hccaef3d5695e586b,64'h40826a44b7edc13f,64'h779eff60c3745b2d,64'h784b4f47d357ef23,
64'hb24afd4a3dfd3e5c,64'hde4aa33b9240e17b,64'hc1fed6b24c0e27d4,64'h4928fd00501ca1d9,
64'h3a62acae5f0a9f5f,64'h56f6f177dffba844,64'h87f11217c5f0ad9b,64'h430b695880d2b06e,
64'h3692662925e33de1,64'h0e25e373023f57d5,64'hbbda236ee22f4bf9,64'hea56ed0a4bb1615e,
64'he9acae8d4aed7994,64'h987633d622722e60,64'h778624a17db43d6e,64'hff7fffff00000081,
64'h003c0cc70d1e41c2,64'h6d978d1c09445e62,64'h2eae706d47a1a370,64'h7bf794dd59d08f8b,
64'h78d5769b6f6a1b00,64'hb520704635472865,64'ha2c6a5a469a038ec,64'hc82e8152e208fa70,
64'h270526cbe222d68d,64'hd5382041476d66a7,64'h4c5c92edd9f1ce34,64'ha6bd70a9fbc19846,
64'h1044b9ce1100dd15,64'h51919d27a229fd65,64'h2640325b803a2278,64'h1f46fe927473c0f8,
64'h649c2623b8ed497f,64'h08e1dd39f4b32822,64'hb6338c7e3f86f116,64'h3811262fc3549f5a,
64'hb80be2f267dcaa9c,64'h06e2a21e937a7623,64'hb0bf717007907c99,64'hf3d91f45685289d2,
64'h73c2d64a53251081,64'h988edf6c8ba5bbc3,64'h7f5bdda8fc98e483,64'h4c56a98e3537dd43,
64'hbe89f1dba58316c8,64'h36e6ee0a706c8023,64'h2490664cb02aed4e,64'h0001fffffffe0000,
64'hae68cf61c7636600,64'h4fcf0b4d85043308,64'h685a3f7a8035a252,64'he57384be5aaf1e77,
64'h9c657fea81ce740f,64'h007bf9646838ea76,64'hf65908fc5b886c79,64'h6aa06f77b298d73f,
64'had9ac9b69653588a,64'h56940147689c9fb2,64'h074fcaa4fbd67572,64'h2deb8ca0773b9aea,
64'h65779eb14af2c352,64'h04135227bf6e09f6,64'hbcf7fb091ba2d965,64'hc25a7a419abf7915,
64'h9257ea56efe9f2db,64'hf25519e292070bd2,64'h0ff6b59860713e9a,64'h4947e80480e50ec6,
64'hd3156573f854faf7,64'hb7b78bc0ffdd421e,64'h3f8890c22f856cd4,64'h185b4ac60695836e,
64'hb493314a2f19ef07,64'h712f1b9811fabea8,64'hded11b7c117a5fc3,64'h52b768595d8b0ae9,
64'h4d657471576bcc99,64'hc3b19eb5139172fc,64'hbc31250eeda1eb6d,64'hfbffffff00000401,
64'h01e0663868f20e10,64'h6cbc68e34a22f30d,64'h7573836b3d0d1b7f,64'hdfbca6edce847c55,
64'hc6abb4de7b50d7fd,64'ha9038236aa394323,64'h16352d284d01c75b,64'h41740a9d1047d37a,
64'h382936601116b467,64'ha9c102103b6b3532,64'h62e49770cf8e719e,64'h35eb8554de0cc22b,
64'h8225ce708806e8a8,64'h8c8ce93f114feb26,64'h320192dd01d113bf,64'hfa37f493a39e07c0,
64'h24e13120c76a4bf5,64'h470ee9cfa5994110,64'hb19c63f6fc3788ab,64'hc089317f1aa4facf,
64'hc05f17983ee554db,64'h371510f49bd3b118,64'h85fb8b853c83e4c3,64'h9ec8fa3242944e89,
64'h9e16b25599288405,64'hc476fb685d2dde14,64'hfadeed4ae4c72415,64'h62b54c73a9beea16,
64'hf44f8ee22c18b63b,64'hb737705483640117,64'h2483326681576a6f,64'h000ffffffff00000,
64'h73467b133b1b2ffb,64'h7e785a6e2821983e,64'h42d1fbd701ad128d,64'h2b9c25f9d578f3b1,
64'he32bff580e73a074,64'h03dfcb2341c753b0,64'hb2c847e9dc4363c1,64'h55037bc094c6b9f5,
64'h6cd64db9b29ac44b,64'hb4a00a3d44e4fd8e,64'h3a7e5527deb3ab90,64'h6f5c6504b9dcd74f,
64'h2bbcf58d57961a8d,64'h209a913dfb704fb0,64'he7bfd84ddd16cb23,64'h12d3d212d5fbc8a2,
64'h92bf52bb7f4f96d4,64'h92a8cf1b90385e89,64'h7fb5acc30389f4d0,64'h4a3f40260728762e,
64'h98ab2ba5c2a7d7b2,64'hbdbc5e0cfeea10eb,64'hfc4486127c2b669f,64'hc2da563034ac1b70,
64'ha4998a5678cf7833,64'h8978dcc38fd5f53d,64'hf688dbe68bd2fe12,64'h95bb42ccec585746,
64'h6b2ba38cbb5e64c6,64'h1d8cf5ae9c8b97da,64'he189287c6d0f5b63,64'hdfffffff00002001,
64'h0f0331c347907080,64'h65e3471d51179865,64'hab9c1b5ce868dbf5,64'hfde537747423e2a2,
64'h355da6f9da86bfe2,64'h481c11ba51ca1913,64'hb1a96942680e3ad8,64'h0ba054ea823e9bce,
64'hc149b30188b5a337,64'h4e081086db59a98b,64'h1724bb897c738ced,64'haf5c2aa7f0661157,
64'h112e73884037453c,64'h646749fc8a7f592c,64'h900c96e90e889df7,64'hd1bfa4a41cf03df9,
64'h270989073b525fa7,64'h38774e7f2cca087e,64'h8ce31fbce1bc4553,64'h04498bfed527d672,
64'h02f8bcc7f72aa6d2,64'hb8a887a5de9d88bf,64'h2fdc5c2de41f2614,64'hf647d19614a27444,
64'hf0b592b0c9442024,64'h23b7db48e96ef09a,64'hd6f76a5e263920a1,64'h15aa63a04df750ad,
64'ha27c771860c5b1d1,64'hb9bb82a91b2008b3,64'h241993350abb5377,64'h007fffffff800000,
64'h9a33d89cd8d97fd5,64'hf3c2d374410cc1ed,64'h168fdeba0d689466,64'h5ce12fcfabc79d87,
64'h195ffac7739d0399,64'h1efe591a0e3a9d80,64'h96423f53e21b1e03,64'ha81bde06a635cfa6,
64'h66b26dd094d62255,64'ha50051ef2727ec6b,64'hd3f2a93ff59d5c7f,64'h7ae32828cee6ba75,
64'h5de7ac6bbcb0d467,64'h04d489f0db827d7f,64'h3dfec275e8b65911,64'h969e9096afde4510,
64'h95fa95dffa7cb69c,64'h954678e081c2f444,64'hfdad661b1c4fa67d,64'h51fa01323943b16e,
64'hc5595d32153ebd8c,64'hede2f06cf7508753,64'he224309ae15b34f1,64'h16d2b187a560db7a,
64'h24cc52b8c67bc193,64'h4bc6e6207eafa9e4,64'hb446df3b5e97f089,64'hadda166b62c2ba2c,
64'h595d1c68daf3262d,64'hec67ad74e45cbed0,64'h0c4943ea687adb11,64'hfffffffe00010002,
64'h78198e1a3c838400,64'h2f1a38ed88bcc325,64'h5ce0daec4346dfa3,64'hef29bbaaa11f1509,
64'haaed37cfd435ff0f,64'h40e08dd48e50c896,64'h8d4b4a184071d6bb,64'h5d02a75411f4de70,
64'h0a4d981245ad19b2,64'h70408438dacd4c56,64'hb925dc4be39c6768,64'h7ae1554483308ab3,
64'h89739c4201ba29e0,64'h233a4fe753fac95d,64'h8064b74c7444efb4,64'h8dfd2526e781efc2,
64'h384c483ada92fd37,64'hc3ba73fa665043ef,64'h6718fdeb0de22a94,64'h224c5ff6a93eb390,
64'h17c5e63fb9553690,64'hc5443d33f4ec45f3,64'h7ee2e17020f9309f,64'hb23e8cb7a513a219,
64'h85ac958d4a210119,64'h1dbeda484b7784cf,64'hb7bb52f731c90502,64'had531d026fba8568,
64'h13e3b8c8062d8e83,64'hcddc154dd9004593,64'h20cc99a955da9bb7,64'h03fffffffc000000,
64'hd19ec4eac6cbfea4,64'h9e169ba908660f61,64'hb47ef5d06b44a330,64'he7097e7f5e3cec36,
64'hcaffd63b9ce81cc8,64'hf7f2c8d071d4ec00,64'hb211faa310d8f014,64'h40def03a31ae7d2b,
64'h35936e87a6b112a5,64'h28028f7e393f6353,64'h9f954a05aceae3f2,64'hd71941497735d3a5,
64'hef3d635fe586a336,64'h26a44f86dc13ebf8,64'heff613b045b2c887,64'hb4f484b97ef2287c,
64'hafd4af03d3e5b4dc,64'haa33c7080e17a21c,64'hed6b30dfe27d33e1,64'h8fd00993ca1d8b6e,
64'h2acae996a9f5ec5a,64'h6f17836eba843a91,64'h112184de0ad9a781,64'hb6958c3d2b06dbd0,
64'h266295c733de0c97,64'h5e373105f57d4f1e,64'ha236f9dff4bf8443,64'h6ed0b3601615d15b,
64'hcae8e348d7993166,64'h633d6bae22e5f679,64'h624a1f5343d6d888,64'hfffffff700080009,
64'hc0cc70d4e41c1ffd,64'h78d1c76d45e61927,64'he706d7641a36fd16,64'h794ddd5c08f8a841,
64'h5769be83a1aff873,64'h07046ea6728644ae,64'h6a5a50c6038eb5d4,64'he8153aa28fa6f37e,
64'h526cc0922d68cd90,64'h820421c9d66a62ad,64'hc92ee2641ce33b3b,64'hd70aaa2719845595,
64'h4b9ce2140dd14efc,64'h19d27f3b9fd64ae7,64'h0325ba67a2277d9c,64'h6fe9293b3c0f7e0c,
64'hc26241d7d497e9b7,64'h1dd39fd932821f72,64'h38c7ef5b6f11549d,64'h1262ffb649f59c7f,
64'hbe2f31fdcaa9b480,64'h2a21e9a5a7622f92,64'hf7170b8407c984f5,64'h91f465c2289d10c3,
64'h2d64ac6e510808c4,64'hedf6d2425bbc2678,64'hbdda97be8e48280b,64'h6a98e8187dd42b3b,
64'h9f1dc640316c7418,64'h6ee0aa74c8022c92,64'h0664cd4baed4ddb7,64'h1fffffffe0000000,
64'h8cf6275c365ff51a,64'hf0b4dd4c43307b04,64'ha3f7ae885a25197b,64'h384bf401f1e761a9,
64'h57feb1e2e740e63a,64'hbf96468a8ea75ff9,64'h908fd51d86c7809b,64'h06f781d38d73e956,
64'hac9b743e35889527,64'h40147bf2c9fb1a97,64'hfcaa503167571f8c,64'hb8ca0a51b9ae9d22,
64'h79eb1b062c3519a9,64'h35227c37e09f5fbf,64'h7fb09d892d964431,64'ha7a425d0f79143db,
64'h7ea578239f2da6db,64'h519e384570bd10db,64'h6b59870613e99f01,64'h7e804ca250ec5b6c,
64'h56574cb64faf62cf,64'h78bc1b78d421d485,64'h890c26f056cd3c08,64'hb4ac61ee5836de7b,
64'h3314ae3a9ef064b7,64'hf1b98831abea78ee,64'h11b7cf04a5fc2213,64'h76859b03b0ae8ad5,
64'h57471a4cbcc98b2a,64'h19eb5d74172fb3c5,64'h1250fa9d1eb6c43d,64'hffffffbf00400041,
64'h066386ad20e0ffe2,64'hc68e3b6d2f30c935,64'h3836bb27d1b7e8a9,64'hca6eeae347c54205,
64'hbb4df41f0d7fc396,64'h3823753394322570,64'h52d286331c75ae9d,64'h40a9d51b7d379be9,
64'h936604936b466c7e,64'h10210e52b3531564,64'h49771326e719d9d2,64'hb855513ecc22aca2,
64'h5ce710a26e8a77de,64'hce93f9dcfeb25738,64'h192dd33d113bece0,64'h7f4949dce07bf05d,
64'h13120ec4a4bf4db2,64'hee9cfec99410fb90,64'hc63f7adc788aa4e7,64'h9317fdb24face3f8,
64'hf1798ff3554da3fb,64'h510f4d2e3b117c8f,64'hb8b85c273e4c27a1,64'h8fa32e1544e88614,
64'h6b2563738840461f,64'h6fb69219dde133b9,64'heed4bdf972414053,64'h54c740c6eea159d5,
64'hf8ee32058b63a0bc,64'h770553a94011648d,64'h33266a5d76a6edb8,64'hffffffff00000000,
64'h67b13ae5b2ffa8cc,64'h85a6ea691983d819,64'h1fbd7447d128cbd3,64'hc25fa0108f3b0d47,
64'hbff58f193a0731ce,64'hfcb23459753affc3,64'h847ea8f0363c04d4,64'h37bc0e9c6b9f4ab0,
64'h64dba1f6ac44a933,64'h00a3df984fd8d4b6,64'he55281923ab8fc59,64'hc6505292cd74e90b,
64'hcf58d83461a8cd45,64'ha913e1c004fafdf7,64'hfd84ec4c6cb22185,64'h3d212e8cbc8a1ed3,
64'hf52bc11ff96d36d5,64'h8cf1c22d85e886d6,64'h5acc38339f4cf805,64'hf40265158762db5d,
64'hb2ba65b47d7b1676,64'hc5e0dbc9a10ea425,64'h48613786b669e03c,64'ha5630f77c1b6f3d3,
64'h98a571d5f78325b7,64'h8dcc41945f53c769,64'h8dbe78252fe11098,64'hb42cd820857456a5,
64'hba38d267e64c594e,64'hcf5aeba0b97d9e28,64'h9287d4e8f5b621e8,64'hfffffdff02000201,
64'h331c35690707ff10,64'h3471db6f798649a2,64'hc1b5d93f8dbf4547,64'h537757203e2a1022,
64'hda6fa0fd6bfe1cab,64'hc11ba99da1912b7f,64'h9694319ae3ad74e6,64'h054ea8dde9bcdf46,
64'h9b30249f5a3363ec,64'h810872959a98ab20,64'h4bb8993938cece8e,64'hc2aa89fb6115650b,
64'he73885157453beee,64'h749fceedf592b9ba,64'hc96e99e889df6700,64'hfa4a4eea03df82e5,
64'h9890762525fa6d90,64'h74e7f653a087dc79,64'h31fbd6e9c4552732,64'h98bfed967d671fbc,
64'h8bcc7fa1aa6d1fd1,64'h887a6973d88be476,64'hc5c2e13ef2613d03,64'h7d1970ae2744309c,
64'h592b1b9f420230f5,64'h7db490d1ef099dc5,64'h76a5efd2920a0291,64'ha63a0639750acea6,
64'hc77190335b1d05d9,64'hb82a9d4d008b2465,64'h993352ecb5376dbf,64'hfffffffefffffff9,
64'h3d89d73097fd465d,64'h2d37534ccc1ec0c4,64'hfdeba23e89465e98,64'h12fd008a79d86a32,
64'hffac78ced0398e6b,64'he591a2d2a9d7fe11,64'h23f54785b1e0269c,64'hbde074e45cfa557f,
64'h26dd0fb862254995,64'h051efcc27ec6a5b0,64'h2a940c98d5c7e2c1,64'h3282949c6ba74852,
64'h7ac6c1a90d466a22,64'h489f0e0527d7efb3,64'hec27626a65910c21,64'he9097466e450f697,
64'ha95e0906cb69b6a1,64'h678e11702f4436ac,64'hd661c19efa67c026,64'ha01328b33b16dae1,
64'h95d32da8ebd8b3ab,64'h2f06de5308752122,64'h4309bc37b34f01de,64'h2b187bc30db79e93,
64'hc52b8eb3bc192db4,64'h6e620ca6fa9e3b44,64'h6df3c12d7f0884bc,64'ha166c1092ba2b523,
64'hd1c693443262ca6b,64'h7ad75d0bcbecf13a,64'h943ea74badb10f3c,64'hffffefff10001001,
64'h98e1ab49383ff87f,64'ha38edb7ccc324d0f,64'h0daeca026dfa2a32,64'h9bbab903f150810e,
64'hd37d07f15ff0e552,64'h08dd4cf30c895bf2,64'hb4a18cdb1d6ba72c,64'h2a7546ef4de6fa30,
64'hd98124fed19b1f5c,64'h084394b0d4c558fc,64'h5dc4c9cbc676746e,64'h15544fe108ab2852,
64'h39c428b2a29df769,64'ha4fe7772ac95cdcd,64'h4b74cf4a4efb37fa,64'hd25277571efc1721,
64'hc483b12d2fd36c7c,64'ha73fb2a0043ee3c5,64'h8fdeb74f22a9398f,64'hc5ff6cb7eb38fddc,
64'h5e63fd115368fe84,64'h43d34ba2c45f23ac,64'h2e1709fd9309e812,64'he8cb85743a2184dd,
64'hc958dcfc101187a6,64'heda48692784cee25,64'hb52f7e9790501485,64'h31d031d0a856752b,
64'h3b8c81a0d8e82ec2,64'hc154ea6d04592323,64'hc99a9769a9bb6df4,64'hfffffffeffffffc1,
64'hec4eb985bfea32e7,64'h69ba9a6760f6061f,64'hef5d11fb4a32f4b9,64'h97e80453cec35190,
64'hfd63c67d81cc7351,64'h2c8d169c4ebff081,64'h1faa3c2e8f0134df,64'hef03a727e7d2abf3,
64'h36e87dc4112a4ca7,64'h28f7e613f6352d80,64'h54a064c7ae3f1607,64'h9414a4e45d3a428f,
64'hd6360d4b6a33510d,64'h44f8702b3ebf7d96,64'h613b135a2c886101,64'h484ba33e2287b4b1,
64'h4af0483b5b4db503,64'h3c708b847a21b55d,64'hb30e0cfdd33e012a,64'h0099459ed8b6d703,
64'hae996d4b5ec59d54,64'h7836f29943a9090f,64'h184de1bf9a780eee,64'h58c3de196dbcf497,
64'h295c75a3e0c96d9a,64'h7310653ad4f1da1d,64'h6f9e096ef84425dd,64'h0b36084e5d15a913,
64'h8e349a2793165352,64'hd6bae8615f6789cd,64'ha1f53a616d8879dc,64'hffff7fff80008001,
64'hc70d5a4dc1ffc3f4,64'h1c76dbeb61926873,64'h6d7650136fd15190,64'hddd5c8238a84086c,
64'h9be83f90ff872a8a,64'h46ea6798644adf90,64'ha50c66ddeb5d395b,64'h53aa377b6f37d17f,
64'hcc0927fc8cd8fada,64'h421ca586a62ac7e0,64'hee264e6033b3a36e,64'haaa27f0845594290,
64'hce21459614efbb47,64'h27f3bb9a64ae6e63,64'h5ba67a5477d9bfce,64'h9293babef7e0b902,
64'h241d896f7e9b63da,64'h39fd950521f71e23,64'h7ef5ba7d1549cc74,64'h2ffb65c559c7eeda,
64'hf31fe88c9b47f41e,64'h1e9a5d1822f91d5e,64'h70b84fed984f408f,64'h465c2ba8d10c26e1,
64'h4ac6e7e6808c3d2a,64'h6d24349ac2677121,64'ha97bf4c18280a423,64'h8e818e8642b3a957,
64'hdc640d07c741760f,64'h0aa7536e22c91912,64'h4cd4bb534ddb6f9a,64'hfffffffefffffe01,
64'h6275cc34ff519731,64'h4dd4d33e07b030f5,64'h7ae88fe15197a5c1,64'hbf4022a2761a8c7c,
64'heb1e33f30e639a81,64'h6468b4e375ff8407,64'hfd51e1747809a6f8,64'h781d39463e955f91,
64'hb743ee2189526537,64'h47bf30a0b1a96bff,64'ha503263f71f8b036,64'ha0a52726e9d21474,
64'hb1b06a61519a8862,64'h27c3815bf5fbecae,64'h09d89ad464430805,64'h425d19f3143da586,
64'h578241dcda6da816,64'he3845c24d10daae7,64'h987067f399f0094b,64'h04ca2cf6c5b6b818,
64'h74cb6a5ff62cea9b,64'hc1b794cd1d484875,64'hc26f0dfcd3c07770,64'hc61ef0cd6de7a4b6,
64'h4ae3ad20064b6ccf,64'h988329d9a78ed0e5,64'h7cf04b7ac2212ee5,64'h59b04272e8ad4898,
64'h71a4d14098b29a8c,64'hb5d74310fb3c4e62,64'h0fa9d3106c43cedb,64'hfffc000300040001,
64'h386ad2740ffe1f9a,64'he3b6df5b0c934398,64'h6bb2809e7e8a8c7d,64'heeae41225420435a,
64'hdf41fc8bfc39544c,64'h37533cc52256fc7e,64'h286336f45ae9cad3,64'h9d51bbdd79be8bf6,
64'h60493fea66c7d6ca,64'h10e52c3731563efe,64'h713273089d9d1b69,64'h5513f8472aca147b,
64'h710a2cb6a77dda32,64'h3f9ddcd425737317,64'hdd33d2a5becdfe6e,64'h949dd5fbbf05c80c,
64'h20ec4b7cf4db1ecf,64'hcfeca82a0fb8f117,64'hf7add3ebaa4e639d,64'h7fdb2e2bce3f76cf,
64'h98ff446bda3fa0e9,64'hf4d2e8c117c8eaf0,64'h85c27f6fc27a0475,64'h32e15d4888613706,
64'h56373f360461e94e,64'h6921a4d9133b8905,64'h4bdfa61114052113,64'h740c7436159d4ab4,
64'he32068443a0bb072,64'h553a9b711648c890,64'h66a5da9c6edb7cce,64'hfffffffefffff001,
64'h13ae61aafa8cb985,64'h6ea699f23d8187a6,64'hd7447f0d8cbd2e05,64'hfa011518b0d463db,
64'h58f19f9f731cd401,64'h2345a71eaffc2035,64'hea8f0baac04d37b9,64'hc0e9ca34f4aafc85,
64'hba1f71114a9329b3,64'h3df985078d4b5ff6,64'h281932008fc581ab,64'h0529393c4e90a39b,
64'h8d83530f8cd4430b,64'h3e1c0ae0afdf656f,64'h4ec4d6a322184028,64'h12e8cf9aa1ed2c2e,
64'hbc120ee8d36d40ae,64'h1c22e12d886d5731,64'hc3833fa0cf804a54,64'h265167b62db5c0c0,
64'ha65b5302b16754d5,64'h0dbca66eea4243a2,64'h13786fec9e03bb7a,64'h30f786716f3d25aa,
64'h571d6902325b6676,64'hc4194ed13c768724,64'he7825bd911097725,64'hcd821399456a44be,
64'h8d268a07c594d45d,64'haeba188cd9e2730b,64'h7d4e9883621e76d8,64'hffe0001f00200001,
64'hc35693a17ff0fccf,64'h1db6fadf649a1cb9,64'h5d9404f6f45463e5,64'h75720919a1021ac9,
64'hfa0fe465e1caa25a,64'hba99e62a12b7e3ef,64'h4319b7a3d74e5697,64'hea8ddeefcdf45fac,
64'h0249ff56363eb64d,64'h872961b98ab1f7f0,64'h89939847ece8db45,64'ha89fc23b5650a3d6,
64'h885165b83beed18d,64'hfceee6a22b9b98b7,64'he99e9533f66ff36a,64'ha4eeafe1f82e405c,
64'h07625be8a6d8f677,64'h7f6541567dc788b2,64'hbd6e9f6452731ce1,64'hfed9716171fbb675,
64'hc7fa2362d1fd0744,64'ha697460fbe475779,64'h2e13fb8213d023a4,64'h970aea454309b82f,
64'hb1b9f9b2230f4a6e,64'h490d26cb99dc4825,64'h5efd308aa0290896,64'ha063a1b3acea559d,
64'h19034228d05d8389,64'ha9d4db8ab246447e,64'h352ed4e676dbe66d,64'hfffffffeffff8001,
64'h9d730d57d465cc28,64'h7534cf94ec0c3d2d,64'hba23f87265e97022,64'hd008a8cc86a31ed1,
64'hc78cfcfd98e6a006,64'h1a2d38f67fe101a7,64'h54785d5d0269bdc1,64'h074e51ada557e422,
64'hd0fb888f54994d93,64'hefcc283d6a5affaf,64'h40c990057e2c0d57,64'h2949c9e274851cd8,
64'h6c1a988066a21854,64'hf0e057067efb2b77,64'h7626b51b10c2013e,64'h97467cd50f696170,
64'he090774b9b6a056b,64'he117096c436ab988,64'h1c19fd0c7c02529a,64'h328b3db26dae05ff,
64'h32da981a8b3aa6a3,64'h6de5337752121d10,64'h9bc37f64f01ddbd0,64'h87bc338c79e92d4f,
64'hb8eb481392db33ae,64'h20ca768fe3b4391a,64'h3c12decf884bb921,64'h6c109cd02b5225ea,
64'h693450422ca6a2e4,64'h75d0c46bcf139853,64'hea74c41e10f3b6bd,64'hff0000ff01000001,
64'h1ab49d11ff87e672,64'hedb7d6fb24d0e5c8,64'heca027b9a2a31f26,64'hab9048d00810d645,
64'hd07f23360e5512c9,64'hd4cf315595bf1f73,64'h18cdbd20ba72b4b6,64'h546ef7856fa2fd59,
64'h124ffab1b1f5b268,64'h394b0dd0558fbf7c,64'h4c9cc2436746da24,64'h44fe11dfb2851eab,
64'h428b2dc5df768c64,64'he77735185cdcc5b1,64'h4cf4a9a6b37f9b49,64'h27757f14c17202db,
64'h3b12df4536c7b3b8,64'hfb2a0ab6ee3c458d,64'heb74fb279398e703,64'hf6cb8b128fddb3a1,
64'h3fd11b1c8fe83a1a,64'h34ba3082f23abbc3,64'h709fdc119e811d1f,64'hb857522e184dc174,
64'h8dcfcd96187a536b,64'h4869365ecee24126,64'hf7e98457014844ae,64'h031d0da26752ace3,
64'hc81a114682ec1c48,64'h4ea6dc5a923223eb,64'ha976a734b6df3367,64'hfffffffefffc0001,
64'heb986ac2a32e613c,64'ha9a67caa6061e965,64'hd11fc3982f4b810b,64'h8045466a3518f682,
64'h3c67e7f2c735002a,64'hd169c7b3ff080d38,64'ha3c2eaea134dee06,64'h3a728d6d2abf2110,
64'h87dc4480a4ca6c92,64'h7e6141f252d7fd71,64'h064c802df1606ab6,64'h4a4e4f14a428e6bf,
64'h60d4c4063510c29d,64'h8702b83af7d95bb1,64'hb135a8db861009ed,64'hba33e6ac7b4b0b7c,
64'h0483ba63db502b51,64'h08b84b691b55cc39,64'he0cfe863e01294d0,64'h9459ed946d702ff7,
64'h96d4c0d559d53517,64'h6f299bbd9090e87d,64'hde1bfb2b80eede7c,64'h3de19c67cf496a74,
64'hc75a40a196d99d6b,64'h0653b4801da1c8cf,64'he096f67d425dc907,64'h6084e6845a912f4d,
64'h49a282146535171d,64'hae862361789cc295,64'h53a620f7879db5e1,64'hf80007ff08000001,
64'hd5a4e88ffc3f3390,64'h6dbeb7e026872e39,64'h65013dd41518f929,64'h5c8246854086b223,
64'h83f919b672a89642,64'ha6798ab2adf8fb92,64'hc66de905d395a5b0,64'ha377bc2d7d17eac6,
64'h927fd58d8fad9340,64'hca586e83ac7dfbdf,64'h64e6121d3a36d11e,64'h27f08eff9428f556,
64'h14596e30fbb4631e,64'h3bb9a8c9e6e62d81,64'h67a54d379bfcda46,64'h3babf8a70b9016d7,
64'hd896fa2ab63d9dbf,64'hd95055be71e22c61,64'h5ba7d9439cc73811,64'hb65c589b7eed9d01,
64'hfe88d8e57f41d0cf,64'ha5d1841891d5de17,64'h84fee08ff408e8f5,64'hc2ba9175c26e0b9b,
64'h6e7e6cb4c3d29b54,64'h4349b2f87712092e,64'hbf4c22bf0a422569,64'h18e86d133a956718,
64'h40d08a3a1760e23a,64'h7536e2d691911f56,64'h4bb539aab6f99b33,64'hfffffffeffe00001,
64'h5cc3561c197309d9,64'h4d33e558030f4b23,64'h88fe1cc77a5c0852,64'h022a3355a8c7b40c,
64'he33f3f9739a8014f,64'h8b4e3da5f84069ba,64'h1e1757559a6f702b,64'hd3946b6a55f9087f,
64'h3ee224092653648c,64'hf30a0f9596bfeb85,64'h3264016f8b0355b0,64'h527278a7214735f6,
64'h06a62034a88614e5,64'h3815c1dbbecadd84,64'h89ad46e130804f63,64'hd19f3568da585bdb,
64'h241dd31eda815a88,64'h45c25b48daae61c8,64'h067f43260094a679,64'ha2cf6ca76b817fb4,
64'hb6a606aecea9a8b4,64'h794cddef848743e5,64'hf0dfd9620776f3da,64'hef0ce33f7a4b539f,
64'h3ad20512b6cceb52,64'h329da400ed0e4678,64'h04b7b3f112ee4831,64'h04273425d4897a65,
64'h4d1410a529a8b8e6,64'h74311b10c4e614a3,64'h9d3107be3cedaf06,64'hc0003fff40000001,
64'had274485e1f99c7a,64'h6df5bf04343971c5,64'h2809eea3a8c7c945,64'he412342c04359116,
64'h1fc8cdb79544b20c,64'h33cc559a6fc7dc8b,64'h336f48349cad2d7a,64'h1bbde170e8bf562b,
64'h93feac707d6c99fc,64'h52c3742363efdef2,64'h273090ecd1b688ed,64'h3f8477fda147aaaf,
64'ha2cb7187dda318f0,64'hddcd465037316c07,64'h3d2a69bfdfe6d22d,64'hdd5fc5395c80b6b7,
64'hc4b7d15bb1ecedf2,64'hca82adf98f116302,64'hdd3eca1ee639c086,64'hb2e2c4e0f76ce803,
64'hf446c732fa0e8671,64'h2e8c20c98eaef0b3,64'h27f70483a04747a4,64'h15d48bb413705cd2,
64'h73f365a91e94da9d,64'h1a4d97c5b890496e,64'hfa6115fd52112b43,64'hc7436899d4ab38c0,
64'h068451d2bb0711ce,64'ha9b716b78c88faad,64'h5da9cd57b7ccd996,64'hfffffffeff000001,
64'he61ab0e2cb984ec6,64'h699f2ac2187a5916,64'h47f0e63fd2e0428c,64'h11519aad463da060,
64'h19f9fcc0cd400a71,64'h5a71ed33c2034dcc,64'hf0babaacd37b8158,64'h9ca35b58afc843f2,
64'hf711204a329b245f,64'h98507cb3b5ff5c21,64'h93200b7d581aad7f,64'h9393c53b0a39afae,
64'h353101a54430a728,64'hc0ae0edef656ec1f,64'h4d6a370d84027b14,64'h8cf9ab4cd2c2ded2,
64'h20ee98f7d40ad43f,64'h2e12da48d5730e3e,64'h33fa193004a533c8,64'h167b65405c0bfd9b,
64'hb530357b754d459b,64'hca66ef7f243a1f25,64'h86fecb173bb79ec9,64'h78671a02d25a9cf1,
64'hd6902896b6675a8f,64'h94ed2008687233bf,64'h25bd9f8897724188,64'h2139a12ea44bd328,
64'h68a0852b4d45c72e,64'ha188d8892730a515,64'he9883df5e76d782c,64'h0002000000000002,
64'h693a24340fcce3cb,64'h6fadf824a1cb8e25,64'h404f751e463e4a27,64'h2091a16721ac88a9,
64'hfe466dbcaa259060,64'h9e62acd47e3ee457,64'h9b7a41a5e5696bcf,64'hddef0b8745fab158,
64'h9ff56387eb64cfdc,64'h961ba11d1f7ef78e,64'h398487678db44767,64'hfc23bfee0a3d5577,
64'h165b8c43ed18c77b,64'hee6a3287b98b6032,64'he9534dffff369167,64'heafe29d0e405b5b2,
64'h25be8ae38f676f8a,64'h54156fd2788b180a,64'he9f650fd31ce042a,64'h9716270cbb674013,
64'ha236399ed0743381,64'h7461064d75778597,64'h3fb8241e023a3d1f,64'haea45da09b82e690,
64'h9f9b2d4bf4a6d4e5,64'hd26cbe2dc4824b70,64'hd308aff190895a11,64'h3a1b44d4a559c5fa,
64'h34228e95d8388e70,64'h4db8b5c16447d563,64'hed4e6abfbe66ccae,64'hfffffffef8000001,
64'h30d5871d5cc27629,64'h4cf95613c3d2c8ad,64'h3f8732009702145e,64'h8a8cd56a31ed0300,
64'hcfcfe6066a005388,64'hd38f69a0101a6e5e,64'h85d5d56d9bdc0ab9,64'he51adac97e421f8c,
64'hb889025894d922f1,64'hc283e5a1affae104,64'h99005beec0d56bf4,64'h9c9e29dc51cd7d6c,
64'ha9880d2b2185393f,64'h057076fdb2b760f2,64'h6b51b86e2013d89e,64'h67cd5a6a9616f68c,
64'h0774c7bfa056a1f7,64'h7096d247ab9871ef,64'h9fd0c98125299e3f,64'hb3db2a02e05fecd8,
64'ha981abe0aa6a2cd3,64'h53377bff21d0f922,64'h37f658bdddbcf644,64'hc338d01992d4e785,
64'hb48144bbb33ad472,64'ha769004743919df4,64'h2decfc45bb920c3f,64'h09cd0976225e993f,
64'h4504295d6a2e396d,64'h0c46c44e398528a3,64'h4c41efb63b6bc159,64'h0010000000000010,
64'h49d121a37e671e55,64'h7d6fc1280e5c7125,64'h027ba8f431f25136,64'h048d0b3a0d644547,
64'hf2336dec512c82f9,64'hf31566a7f1f722b4,64'hdbd20d332b4b5e74,64'hef785c402fd58aba,
64'hffab1c435b267edc,64'hb0dd08ecfbf7bc6c,64'hcc243b3d6da23b37,64'he11dff7751eaabb1,
64'hb2dc621f68c63bd8,64'h73519444cc5b0189,64'h4a9a7006f9b48b31,64'h57f14e8e202dad89,
64'h2df4571d7b3b7c4f,64'ha0ab7e95c458c04e,64'h4fb287f08e702149,64'hb8b13869db3a0094,
64'h11b1ccfb83a19c03,64'ha308326eabbc2cb5,64'hfdc120f111d1e8f7,64'h7522ed09dc17347b,
64'hfcd96a63a536a724,64'h9365f17424125b7a,64'h98457f92844ad082,64'hd0da26a62ace2fcf,
64'ha11474afc1c4737f,64'h6dc5ae0d223eab16,64'h6a735604f3366569,64'hfffffffec0000001,
64'h86ac38ebe613b147,64'h67cab0a01e964566,64'hfc399005b810a2ef,64'h5466ab558f6817fc,
64'h7e7f303950029c3a,64'h9c7b4d0680d372ea,64'h2eaeab70dee055c4,64'h28d6d652f210fc59,
64'hc44812c9a6c91783,64'h141f2d137fd7081a,64'hc802df7a06ab5f9c,64'he4f14ee68e6beb5c,
64'h4c40695e0c29c9f3,64'h2b83b7ed95bb0790,64'h5a8dc374009ec4ed,64'h3e6ad357b0b7b45d,
64'h3ba63dfd02b50fb8,64'h84b692405cc38f75,64'hfe864c0d294cf1f4,64'h9ed9501c02ff66bb,
64'h4c0d5f0a53516693,64'h99bbdffb0e87c90e,64'hbfb2c5efede7b21f,64'h19c680d296a73c22,
64'ha40a25e299d6a38b,64'h3b48023f1c8cef9b,64'h6f67e22edc9061f7,64'h4e684bb112f4c9f8,
64'h28214aed5171cb66,64'h62362271cc294518,64'h620f7db3db5e0ac6,64'h0080000000000080,
64'h4e890d1df338f2a6,64'heb7e094372e38925,64'h13dd47a18f9289b0,64'h246859d06b222a38,
64'h919b6f69896417c1,64'h98ab35468fb91599,64'hde90699f5a5af39a,64'h7bc2e2087eac55c9,
64'hfd58e221d933f6d9,64'h86e8476cdfbde35b,64'h6121d9f16d11d9b2,64'h08effbc18f555d81,
64'h96e311004631debb,64'h9a8ca22962d80c45,64'h54d38039cda45986,64'hbf8a7473016d6c46,
64'h6fa2b8ecd9dbe277,64'h055bf4b322c6026b,64'h7d943f8673810a46,64'hc589c353d9d0049b,
64'h8d8e67dc1d0ce018,64'h1841937a5de165a3,64'hee09078f8e8f47b1,64'ha9176851e0b9a3d5,
64'he6cb532429b53919,64'h9b2f8ba52092dbcc,64'hc22bfc982256840c,64'h86d1353756717e72,
64'h08a3a5830e239bf3,64'h6e2d706c11f558ad,64'h539ab02a99b32b45,64'hfffffffd00000001,
64'h3561c763309d8a34,64'h3e558503f4b22b2d,64'he1cc8034c0851771,64'ha3355aae7b40bfde,
64'hf3f981cd8014e1cd,64'he3da6838069b974c,64'h75755b87f702ae1f,64'h46b6b2989087e2c7,
64'h224096533648bc12,64'ha0f9689bfeb840d0,64'h4016fbd6355afcda,64'h278a773b735f5ad9,
64'h62034af2614e4f96,64'h5c1dbf6dadd83c7f,64'hd46e1ba204f62766,64'hf3569abe85bda2e7,
64'hdd31efe915a87dbf,64'h25b49206e61c7ba4,64'hf43260704a678f99,64'hf6ca80e417fb35d4,
64'h606af8549a8b3496,64'hcddeffdc743e486c,64'hfd962f846f3d90f3,64'hce340694b539e110,
64'h20512f19ceb51c53,64'hda4011f9e4677cd7,64'h7b3f1179e4830fb5,64'h73425d8a97a64fbe,
64'h410a576b8b8e5b2f,64'h11b11391614a28bd,64'h107beda1daf0562d,64'h0400000000000400,
64'h744868f199c7952e,64'h5bf04a22971c4921,64'h9eea3d0c7c944d80,64'h2342ce84591151bf,
64'h8cdb7b504b20be04,64'hc559aa387dc8acc4,64'hf4834d00d2d79cca,64'hde171046f562ae45,
64'heac71115c99fb6c1,64'h37423b6afdef1ad4,64'h090ecf8e688ecd8d,64'h477fde0c7aaaec08,
64'hb7188806318ef5d4,64'hd465114f16c06224,64'ha69c01d06d22cc2e,64'hfc53a39d0b6b622b,
64'h7d15c769cedf13b5,64'h2adfa59916301358,64'heca1fc369c08522d,64'h2c4e1aa4ce8024d2,
64'h6c733ee4e86700bc,64'hc20c9bd2ef0b2d18,64'h70483c83747a3d81,64'h48bb429405cd1ea3,
64'h365a99284da9c8c1,64'hd97c5d2d0496de5c,64'h115fe4c712b4205a,64'h3689a9beb38bf38c,
64'h451d2c18711cdf98,64'h716b83638faac565,64'h9cd58156cd995a26,64'hffffffef00000001,
64'hab0e3b1a84ec519f,64'hf2ac2820a5915967,64'h0e6401ad0428bb81,64'h19aad578da05feeb,
64'h9fcc0e7300a70e61,64'h1ed341c734dcba59,64'habaadc42b81570f5,64'h35b594c6843f1636,
64'h1204b29ab245e08f,64'h07cb44e4f5c2067b,64'h00b7deb3aad7e6ce,64'h3c53b9dc9afad6c7,
64'h101a57960a727cad,64'he0edfb6f6ec1e3f6,64'ha370dd1627b13b2a,64'h9ab4d5fb2ded1731,
64'he98f7f4ead43edf2,64'h2da4903830e3dd1f,64'ha1930389533c7cc1,64'hb6540727bfd9ae99,
64'h0357c2a7d459a4ad,64'h6ef7fee9a1f2435a,64'hecb17c2a79ec8791,64'h71a034aba9cf087a,
64'h028978cf75a8e297,64'hd2008fd5233be6b2,64'hd9f88bd224187da5,64'h9a12ec57bd327ded,
64'h0852bb5e5c72d976,64'h8d889c8b0a5145e8,64'h83df6d0ed782b168,64'h2000000000002000,
64'ha243478fce3ca96d,64'hdf825116b8e24906,64'hf751e867e4a26bfc,64'h1a167423c88a8df7,
64'h66dbda865905f01c,64'h2acd51c9ee45661a,64'ha41a680d96bce649,64'hf0b8823dab157222,
64'h563888b54cfdb601,64'hba11db58ef78d69f,64'h48767c7344766c68,64'h3bfef065d557603e,
64'hb8c440368c77ae9b,64'ha3288a7eb603111a,64'h34e00e886916616b,64'he29d1cef5b5b1151,
64'he8ae3b5176f89da5,64'h56fd2cc9b1809abf,64'h650fe1bbe0429161,64'h6270d5277401268f,
64'h6399f72a433805dd,64'h1064de9d785968ba,64'h8241e41ea3d1ec05,64'h45da14a22e68f516,
64'hb2d4c9436d4e4607,64'hcbe2e96e24b6f2da,64'h8aff263895a102d0,64'hb44d4df69c5f9c5f,
64'h28e960c588e6fcbe,64'h8b5c1b1f7d562b25,64'he6ac0aba6ccad12c,64'hffffff7f00000001,
64'h5871d8d927628cf3,64'h9561410c2c8acb31,64'h73200d682145dc08,64'hcd56abc6d02ff758,
64'hfe60739c05387304,64'hf69a0e39a6e5d2c8,64'h5d56e21ac0ab87a3,64'hadaca63521f8b1af,
64'h902594d5922f0478,64'h3e5a2727ae1033d8,64'h05bef59d56bf3670,64'he29dcee5d7d6b637,
64'h80d2bcb05393e568,64'h076fdb82760f1fa9,64'h1b86e8b63d89d94b,64'hd5a6afdd6f68b984,
64'h4c7bfa7c6a1f6f89,64'h6d2481c2871ee8f7,64'h0c981c4f99e3e603,64'hb2a03942fecd74c3,
64'h1abe153ea2cd2568,64'h77bff7500f921acd,64'h658be15acf643c81,64'h8d01a5604e7843cd,
64'h144bc67bad4714b8,64'h90047eaf19df358a,64'hcfc45e9720c3ed22,64'hd09762c1e993ef64,
64'h4295daf2e396cbb0,64'h6c44e45c528a2f3c,64'h1efb687abc158b3c,64'h000000010000ffff,
64'h121a3c8371e54b63,64'hfc1288bbc712482a,64'hba8f434625135fd9,64'hd0b3a11e44546fb8,
64'h36ded435c82f80dd,64'h566a8e50722b30cf,64'h20d34071b5e73243,64'h85c411f458ab9109,
64'hb1c445ac67edb006,64'hd08edacc7bc6b4f3,64'h43b3e39c23b3633e,64'hdff7832faabb01ef,
64'hc62201b963bd74d3,64'h194453fab01888cb,64'ha700744448b30b57,64'h14e8e781dad88a81,
64'h4571da92b7c4ed21,64'hb7e9664f8c04d5f6,64'h287f0de202148b05,64'h1386a93ea0093475,
64'h1ccfb95519c02ee5,64'h8326f4ebc2cb45d0,64'h120f20f91e8f6024,64'h2ed0a5137347a8ae,
64'h96a64a206a723033,64'h5f174b7725b796ca,64'h57f931c8ad08167c,64'ha26a6fb9e2fce2f3,
64'h474b062d4737e5ef,64'h5ae0d8ffeab15924,64'h356055da66568959,64'hfffffbff00000001,
64'hc38ec6cb3b146796,64'hab0a086564565984,64'h99006b440a2ee03d,64'h6ab55e3c817fbaba,
64'hf3039ce729c39819,64'hb4d071d4372e9639,64'heab710d8055c3d16,64'h6d6531ae0fc58d73,
64'h812ca6b0917823bc,64'hf2d1393e70819ebf,64'h2df7aceab5f9b380,64'h14ee7735beb5b1b1,
64'h0695e5869c9f2b3c,64'h3b7edc13b078fd48,64'hdc3745b1ec4eca58,64'had357ef17b45cc1a,
64'h63dfd3e550fb7c46,64'h69240e1738f747b5,64'h64c0e27ccf1f3018,64'h9501ca1cf66ba613,
64'hd5f0a9f516692b40,64'hbdffba837c90d665,64'h2c5f0ad97b21e405,64'h680d2b0673c21e64,
64'ha25e33dd6a38a5c0,64'h8023f57ccef9ac4c,64'h7e22f4bf061f690a,64'h84bb16154c9f7b1a,
64'h14aed7991cb65d7e,64'h622722e5945179dd,64'hf7db43d5e0ac59e0,64'h000000080007fff8,
64'h90d1e41b8f2a5b18,64'he09445e538924149,64'hd47a1a36289afec3,64'h859d08f822a37dba,
64'hb6f6a1af417c06e7,64'hb354728591598676,64'h069a038eaf399217,64'h2e208fa6c55c8844,
64'h8e222d683f6d802b,64'h8476d669de35a792,64'h1d9f1ce31d9b19ee,64'hffbc198355d80f72,
64'h31100dd11deba692,64'hca229fd580c44658,64'h3803a22745985ab3,64'ha7473c0ed6c45408,
64'h2b8ed497be276906,64'hbf4b32816026afab,64'h43f86f1110a45827,64'h9c3549f50049a3a8,
64'he67dcaa8ce017728,64'h1937a762165a2e7c,64'h907907c8f47b0120,64'h7685289c9a3d456f,
64'hb532510753918194,64'hf8ba5bbb2dbcb64e,64'hbfc98e476840b3de,64'h13537dd417e71793,
64'h3a58316c39bf2f76,64'hd706c801558ac91e,64'hab02aed432b44ac7,64'hffffdfff00000001,
64'h1c76365fd8a33caa,64'h5850433022b2cc1b,64'hc8035a24517701e4,64'h55aaf1e70bfdd5cd,
64'h981ce7404e1cc0c1,64'ha6838ea6b974b1c3,64'h55b886c72ae1e8a9,64'h6b298d737e2c6b95,
64'h096535888bc11ddc,64'h9689c9fa840cf5f1,64'h6fbd6756afcd9bff,64'ha773b9adf5ad8d88,
64'h34af2c34e4f959e0,64'hdbf6e09e83c7ea3f,64'he1ba2d95627652ba,64'h69abf790da2e60cb,
64'h1efe9f2d87dbe22d,64'h492070bcc7ba3da5,64'h260713e978f980bd,64'ha80e50ebb35d3094,
64'haf854faeb34959fa,64'heffdd420e486b323,64'h62f856ccd90f2027,64'h406958369e10f31d,
64'h12f19ef051c52dfb,64'h011fabea77cd625c,64'hf117a5fb30fb484d,64'h25d8b0ae64fbd8cc,
64'ha576bcc8e5b2ebf0,64'h1139172fa28bcee5,64'hbeda1eb60562cef9,64'h00000040003fffc0,
64'h868f20e07952d8bc,64'h04a22f30c4920a41,64'ha3d0d1b744d7f612,64'h2ce847c5151bedcc,
64'hb7b50d7f0be03733,64'h9aa394318acc33ab,64'h34d01c7579cc90b8,64'h71047d372ae4421f,
64'h71116b45fb6c0154,64'h23b6b352f1ad3c8c,64'hecf8e718ecd8cf70,64'hfde0cc21aec07b89,
64'h88806e89ef5d348f,64'h5114feb2062232ba,64'hc01d113b2cc2d597,64'h3a39e07bb622a03b,
64'h5c76a4bef13b482f,64'hfa59941001357d53,64'h1fc3788a8522c136,64'he1aa4fac024d1d3c,
64'h33ee554d700bb939,64'hc9bd3b10b2d173e0,64'h83c83e4ba3d808fc,64'hb42944e7d1ea2b75,
64'ha992883f9c8c0c9b,64'hc5d2dde06de5b269,64'hfe4c724042059eeb,64'h9a9beea0bf38bc98,
64'hd2c18b62cdf97baf,64'hb8364010ac5648ea,64'h581576a695a25633,64'hfffeffff00000001,
64'he3b1b2fec519e550,64'hc2821983159660d6,64'h401ad1288bb80f1a,64'had578f3a5feeae66,
64'hc0e73a0670e60604,64'h341c753acba58e13,64'hadc4363b570f4546,64'h594c6b9ef1635ca5,
64'h4b29ac445e08eee0,64'hb44e4fd82067af84,64'h7deb3ab87e6cdff5,64'h3b9dcd74ad6c6c3b,
64'ha57961a827caceff,64'hdfb704fa1e3f51f2,64'h0dd16cb213b295c9,64'h4d5fbc89d1730655,
64'hf7f4f96c3edf1168,64'h490385e83dd1ed26,64'h30389f4cc7cc05e7,64'h407287629ae9849b,
64'h7c2a7d7a9a4acfcb,64'h7feea10e24359911,64'h17c2b669c8790135,64'h034ac1b6f08798e6,
64'h978cf7828e296fd8,64'h08fd5f53be6b12e0,64'h88bd2fe087da4261,64'h2ec5857427dec65f,
64'h2bb5e64c2d975f7b,64'h89c8b97d145e7728,64'hf6d0f5b52b1677c3,64'h0000020001fffe00,
64'h34790707ca96c5dc,64'h2511798624905208,64'h1e868dbf26bfb08b,64'h67423e29a8df6e5f,
64'hbda86bfd5f01b993,64'hd51ca19056619d54,64'ha680e3acce6485bf,64'h8823e9bc572210f5,
64'h888b5a32db600a9d,64'h1db59a988d69e45f,64'h67c738ce66c67b79,64'hef0661147603dc41,
64'h440374537ae9a474,64'h88a7f592311195ce,64'h00e889df6616acb2,64'hd1cf03deb11501d7,
64'he3b525f989da4176,64'hd2cca08709abea91,64'hfe1bc454291609b0,64'h0d527d671268e9d9,
64'h9f72aa6c805dc9c7,64'h4de9d88b968b9efa,64'h1e41f2611ec047dc,64'ha14a27438f515ba3,
64'h4c944201e46064d3,64'h2e96ef096f2d9342,64'hf2639209102cf751,64'hd4df7509f9c5e4bc,
64'h960c5b1c6fcbdd72,64'hc1b2008a62b2474b,64'hc0abb536ad12b196,64'hfff7ffff00000001,
64'h1d8d97fd28cf2a79,64'h1410cc1eacb306aa,64'h00d689465dc078ce,64'h6abc79d7ff75732b,
64'h0739d0398730301a,64'ha0e3a9d75d2c7097,64'h6e21b1dfb87a2a2b,64'hca635cf98b1ae526,
64'h594d6224f04776fe,64'ha2727ec6033d7c1b,64'hef59d5c6f366ffa5,64'hdcee6ba66b6361d7,
64'h2bcb0d463e5677f3,64'hfdb827d6f1fa8f8a,64'h6e8b65909d94ae48,64'h6afde4508b9832a6,
64'hbfa7cb68f6f88b39,64'h481c2f43ee8f692e,64'h81c4fa673e602f37,64'h03943b16d74c24d6,
64'he153ebd7d2567e55,64'hff75087421acc885,64'hbe15b34e43c809a8,64'h1a560db7843cc730,
64'hbc67bc18714b7ebc,64'h47eafa9df3589700,64'h45e97f083ed21304,64'h762c2ba23ef632f7,
64'h5daf32626cbafbd7,64'h4e45cbeca2f3b93c,64'hb687adb058b3be11,64'h000010000ffff000,
64'ha3c8383f54b62edf,64'h288bcc322482903f,64'hf4346df935fd8458,64'h3a11f15046fb72f5,
64'hed435feff80dcc93,64'ha8e50c88b30cea9a,64'h34071d6b73242df3,64'h411f4de6b91087a4,
64'h445ad19adb0054e4,64'hedacd4c46b4f22f8,64'h3e39c6763633dbc5,64'h783308aab01ee201,
64'h201ba29dd74d239e,64'h453fac95888cae6c,64'h07444efb30b56590,64'h8e781efb88a80eb2,
64'h1da92fd34ed20ba9,64'h9665043e4d5f5482,64'hf0de22a848b04d79,64'h6a93eb3893474ec8,
64'hfb95536802ee4e34,64'h6f4ec45eb45cf7ce,64'hf20f9308f6023ee0,64'h0a513a217a8add13,
64'h64a2101123032696,64'h74b7784c796c9a0f,64'h931c904f8167ba81,64'ha6fba855ce2f25da,
64'hb062d8e77e5eeb8c,64'h0d90045915923a52,64'h055da9bb68958caa,64'hffbfffff00000001,
64'hec6cbfe9467953c8,64'ha08660f565983550,64'h06b44a32ee03c670,64'h55e3cec2fbab9955,
64'h39ce81cc398180d0,64'h071d4ebfe96384b3,64'h710d8f00c3d15155,64'h531ae7d258d7292a,
64'hca6b1129823bb7ee,64'h1393f63519ebe0d3,64'h7aceae3e9b37fd21,64'he7735d395b1b0eb2,
64'h5e586a32f2b3bf97,64'hedc13ebe8fd47c49,64'h745b2c87eca5723d,64'h57ef22875cc1952d,
64'hfd3e5b4cb7c459c3,64'h40e17a21747b496e,64'h0e27d33df30179b4,64'h1ca1d8b6ba6126b0,
64'h0a9f5ec592b3f2a1,64'hfba843a80d664421,64'hf0ad9a771e404d3b,64'hd2b06dbc21e63980,
64'he33de0c88a5bf5db,64'h3f57d4f19ac4b7fe,64'h2f4bf843f690981e,64'hb1615d14f7b197b5,
64'hed79931565d7deb6,64'h722e5f67179dc9de,64'hb43d6d87c59df083,64'h000080007fff8000,
64'h1e41c1ffa5b176f3,64'h445e6192241481f7,64'ha1a36fd0afec22b9,64'hd08f8a8337db97a7,
64'h6a1aff86c06e6491,64'h4728644a986754cb,64'ha038eb5c99216f97,64'h08fa6f37c8843d1e,
64'h22d68cd8d802a71e,64'h6d66a62a5a7917b9,64'hf1ce33b2b19ede27,64'hc198455880f71005,
64'h00dd14efba691cef,64'h29fd64ae4465735e,64'h3a2277d985ab2c80,64'h73c0f7e04540758c,
64'hed497e9a76905d48,64'hb32821f66afaa40c,64'h86f1154945826bc1,64'h549f59c79a3a763d,
64'hdcaa9b4717727199,64'h7a7622f8a2e7be6d,64'h907c984eb011f6f9,64'h5289d10bd456e898,
64'h2510808c181934ad,64'ha5bbc266cb64d075,64'h98e482800b3dd404,64'h37dd42b371792ecb,
64'h8316c740f2f75c5b,64'h6c8022c8ac91d290,64'h2aed4ddb44ac6550,64'hfdffffff00000001,
64'h6365ff5133ca9e39,64'h043307b02cc1aa7b,64'h35a25197701e3380,64'haf1e7619dd5ccaa6,
64'hce740e62cc0c067f,64'h38ea75ff4b1c2598,64'h886c78091e8a8aa5,64'h98d73e94c6b9494e,
64'h5358895211ddbf6a,64'h9c9fb1a8cf5f0698,64'hd67571f7d9bfe905,64'h3b9ae9d1d8d87589,
64'hf2c35199959dfcb6,64'h6e09f5fb7ea3e241,64'ha2d96442652b91e5,64'hbf79143ce60ca966,
64'he9f2da6cbe22ce11,64'h070bd10da3da4b6e,64'h713e99ef980bcda0,64'he50ec5b5d3093580,
64'h54faf62c959f9508,64'hdd421d476b322101,64'h856cd3bff20269d1,64'h95836de70f31cbfa,
64'h19ef064b52dfaed1,64'hfabea78dd625bfef,64'h7a5fc220b484c0ef,64'h8b0ae8acbd8cbda3,
64'h6bcc98b22ebef5a9,64'h9172fb3bbcee4eed,64'ha1eb6c432cef8413,64'h00040003fffc0000,
64'hf20e0ffd2d8bb798,64'h22f30c9320a40fb6,64'h0d1b7e8a7f6115c3,64'h847c541fbedcbd32,
64'h50d7fc3903732485,64'h39432256c33aa656,64'h01c75ae9c90b7cb3,64'h47d379be4421e8f0,
64'h16b466c7c01538ef,64'h6b353155d3c8bdc5,64'h8e719d9c8cf6f131,64'h0cc22aca07b88022,
64'h06e8a77dd348e778,64'h4feb2573232b9aef,64'hd113becd2d5963ff,64'h9e07bf052a03ac5d,
64'h6a4bf4dab482ea39,64'h99410fb857d5205b,64'h3788aa4e2c135e04,64'ha4face3ed1d3b1e6,
64'he554da3ebb938cc2,64'hd3b117c8173df365,64'h83e4c279808fb7c4,64'h944e8860a2b744be,
64'h28840461c0c9a567,64'h2dde133b5b2683a3,64'hc724140459eea01c,64'hbeea159c8bc97657,
64'h18b63a0b97bae2d4,64'h64011648648e947d,64'h576a6edb25632a7f,64'hefffffff00000001,
64'h1b2ffa8c9e54f1c5,64'h21983d81660d53d8,64'had128cbc80f19bff,64'h78f3b0d3eae6552b,
64'h73a0731c606033f2,64'hc753affb58e12cbf,64'h4363c04cf4545524,64'hc6b9f4aa35ca4a6c,
64'h9ac44a928eedfb4e,64'he4fd8d4a7af834bc,64'hb3ab8fc4cdff4822,64'hdcd74e8fc6c3ac47,
64'h961a8cd3acefe5a9,64'h704fafdef51f1205,64'h16cb2218295c8f23,64'hfbc8a1ec30654b2b,
64'h4f96d36cf1167081,64'h385e886d1ed25b70,64'h89f4cf7fc05e6cfd,64'h28762db59849abf9,
64'ha7d7b166acfca83e,64'hea10ea4159910802,64'h2b669e0390134e84,64'hac1b6f3c798e5fcc,
64'hcf78325a96fd7688,64'hd5f53c75b12dff71,64'hd2fe1108a4260775,64'h58574569ec65ed14,
64'h5e64c59475f7ad45,64'h8b97d9e1e7727764,64'h0f5b621e677c2093,64'h0020001fffe00000,
64'h90707ff06c5dbcb9,64'h1798649a05207daf,64'h68dbf453fb08ae18,64'h23e2a101f6e5e98c,
64'h86bfe1ca1b992426,64'hca1912b719d532af,64'h0e3ad74e485be598,64'h3e9bcdf4210f477e,
64'hb5a3363e00a9c778,64'h59a98ab19e45ee25,64'h738cece867b78984,64'h661156503dc40110,
64'h37453bee9a473bc0,64'h7f592b9b195cd776,64'h889df66f6acb1ff2,64'hf03df82d501d62e4,
64'h525fa6d8a41751c5,64'hca087dc6bea902d4,64'hbc455272609af01f,64'h27d671fb8e9d8f2b,
64'h2aa6d1fcdc9c6609,64'h9d88be46b9ef9b22,64'h1f2613d0047dbe1c,64'ha274430915ba25ec,
64'h4420230f064d2b37,64'h6ef099dbd9341d17,64'h3920a028cf7500da,64'hf750ace95e4bb2b3,
64'hc5b1d05cbdd716a0,64'h2008b2462474a3e5,64'hbb5376db2b1953f6,64'h7fffffff00000001,
64'hd97fd464f2a78e28,64'h0cc1ec0c306a9ebf,64'h689465e9078cdff3,64'hc79d86a25732a955,
64'h9d0398e603019f8d,64'h3a9d7fe0c70965f2,64'h1b1e0269a2a2a91e,64'h35cfa557ae52535a,
64'hd6225498776fda6c,64'h27ec6a5ad7c1a5d9,64'h9d5c7e2b6ffa410b,64'he6ba7484361d6232,
64'hb0d466a1677f2d44,64'h827d7efaa8f89025,64'hb65910c14ae47918,64'hde450f68832a5951,
64'h7cb69b6988b38406,64'hc2f44369f692db7f,64'h4fa67c0202f367e4,64'h43b16dadc24d5fc7,
64'h3ebd8b3a67e541eb,64'h50875211cc884009,64'h5b34f01d809a741f,64'h60db79e8cc72fe5b,
64'h7bc192dab7ebb43a,64'hafa9e3b3896ffb82,64'h97f0884b21303ba2,64'hc2ba2b51632f689e,
64'hf3262ca5afbd6a26,64'h5cbecf133b93bb1c,64'h7adb10f33be10498,64'h010000ffff000000,
64'h8383ff8762ede5c4,64'hbcc324d02903ed78,64'h46dfa2a2d84570bd,64'h1f150810b72f4c5f,
64'h35ff0e54dcc9212c,64'h50c895becea99572,64'h71d6ba7242df2cc0,64'hf4de6fa2087a3bef,
64'had19b1f5054e3bbb,64'hcd4c558ef22f7126,64'h9c6767463dbc4c1d,64'h308ab284ee20087d,
64'hba29df75d239ddff,64'hfac95cdbcae6bbad,64'h44efb37f5658ff8c,64'h81efc17180eb1719,
64'h92fd36c720ba8e26,64'h5043ee3bf548169a,64'he22a939804d780f3,64'h3eb38fdd74ec7957,
64'h55368fe7e4e33047,64'hec45f239cf7cd90c,64'hf9309e8023edf0e0,64'h13a2184dadd12f5b,
64'h2101187a326959b6,64'h7784cee1c9a0e8b5,64'hc90501477ba806cf,64'hba856751f25d9591,
64'h2d8e82ebeeb8b4fa,64'h0045923223a51f27,64'hda9bb6de58ca9fab,64'hfffffffb00000005,
64'hcbfea32d953c713a,64'h660f60618354f5f8,64'h44a32f4b3c66ff95,64'h3cec3518b9954aa2,
64'he81cc734180cfc64,64'hd4ebff07384b2f8f,64'hd8f0134d151548f0,64'hae7d2abe72929acf,
64'hb112a4c9bb7ed35a,64'h3f6352d7be0d2ec7,64'heae3f15f7fd20854,64'h35d3a428b0eb1189,
64'h86a335103bf96a1b,64'h13ebf7d947c48124,64'hb2c8860f5723c8bb,64'hf2287b4a1952ca82,
64'he5b4db4f459c202d,64'h17a21b55b496dbf2,64'h7d33e012179b3f1e,64'h1d8b6d70126afe36,
64'hf5ec59d43f2a0f57,64'h843a909064420046,64'hd9a780ee04d3a0f6,64'h06dbcf496397f2d5,
64'hde0c96d8bf5da1cd,64'h7d4f1da14b7fdc0b,64'hbf84425d0981dd0c,64'h15d15a91197b44ea,
64'h993165347deb5129,64'he5f6789bdc9dd8de,64'hd6d8879cdf0824bd,64'h080007fff8000000,
64'h1c1ffc3f176f2e1c,64'he6192686481f6bbb,64'h36fd1518c22b85e6,64'hf8a84085b97a62f8,
64'haff872a7e649095f,64'h8644adf8754cab8e,64'h8eb5d39516f965fd,64'ha6f37d1743d1df71,
64'h68cd8fad2a71ddd3,64'h6a62ac7d917b892a,64'he33b3a35ede260e4,64'h84559428710043e7,
64'hd14efbb391ceeff3,64'hd64ae6e55735dd61,64'h277d9bfcb2c7fc5e,64'h0f7e0b900758b8c4,
64'h97e9b63d05d4712c,64'h821f71e1aa40b4ce,64'h11549cc726bc0791,64'hf59c7eeca763cab7,
64'ha9b47f4127198236,64'h622f91d57be6c859,64'hc984f4081f6f86f9,64'h9d10c26d6e897ad8,
64'h0808c3d2934acdaf,64'hbc2677114d0745a5,64'h48280a41dd403672,64'hd42b3a9492ecac83,
64'h6c74176075c5a7cf,64'h022c91911d28f938,64'hd4ddb6f8c654fd52,64'hffffffdf00000021,
64'h5ff51972a9e389ca,64'h307b030f1aa7afbd,64'h25197a5be337fca6,64'he761a8c6ccaa550f,
64'h40e639a7c067e319,64'ha75ff83fc2597c72,64'hc7809a6ea8aa477a,64'h73e955f89494d673,
64'h88952652dbf69acb,64'hfb1a96bef0697637,64'h571f8b02fe904299,64'hae9d214687588c47,
64'h3519a885dfcb50d4,64'h9f5fbeca3e240920,64'h9644307fb91e45d3,64'h9143da57ca965409,
64'h2da6da812ce10161,64'hbd10daada4b6df90,64'he99f0093bcd9f8ed,64'hec5b6b809357f1b0,
64'haf62cea8f9507ab1,64'h21d484872210022c,64'hcd3c0776269d07aa,64'h36de7a4b1cbf96a8,
64'hf064b6cbfaed0e62,64'hea78ed0d5bfee055,64'hfc2212ed4c0ee85b,64'hae8ad488cbda2750,
64'hc98b29a7ef5a8944,64'h2fb3c4e5e4eec6e9,64'hb6c43cecf84125e2,64'h40003fffc0000000,
64'he0ffe1f8bb7970e0,64'h30c9343940fb5dd1,64'hb7e8a8c7115c2f2f,64'hc5420434cbd317b9,
64'h7fc3954432484af3,64'h32256fc7aa655c6c,64'h75ae9cacb7cb2fe4,64'h379be8bf1e8efb83,
64'h466c7d6c538eee95,64'h531563ef8bdc494d,64'h19d9d1b66f130719,64'h22aca14788021f34,
64'h8a77dda28e777f92,64'hb2573730b9aeeb02,64'h3becdfe6963fe2ef,64'h7bf05c803ac5c620,
64'hbf4db1ec2ea3895c,64'h10fb8f115205a66c,64'h8aa4e63935e03c88,64'hace3f76c3b1e55b1,
64'h4da3fa0e38cc11ab,64'h117c8eaedf3642c5,64'h4c27a046fb7c37c2,64'he886136f744bd6bc,
64'h40461e949a566d78,64'he133b88f683a2d23,64'h41405210ea01b38e,64'ha159d4aa97656412,
64'h63a0bb06ae2d3e75,64'h11648c88e947c9c0,64'ha6edb7cc32a7ea8a,64'hfffffeff00000101,
64'hffa8cb974f1c4e4e,64'h83d81879d53d7de7,64'h28cbd2e019bfe52f,64'h3b0d463d6552a871,
64'h0731cd40033f18c6,64'h3affc20312cbe38b,64'h3c04d37b45523bca,64'h9f4aafc7a4a6b395,
64'h44a9329adfb4d654,64'hd8d4b5fe834bb1b1,64'hb8fc5819f48214c6,64'h74e90a393ac46233,
64'ha8cd442ffe5a869f,64'hfafdf655f12048fc,64'hb2218401c8f22e94,64'h8a1ed2c254b2a044,
64'h6d36d40a67080b07,64'he886d57225b6fc7b,64'h4cf804a4e6cfc761,64'h62db5c0b9abf8d79,
64'h7b16754cca83d583,64'h0ea4243a1080115f,64'h69e03bb734e83d4a,64'hb6f3d259e5fcb53f,
64'h8325b666d7687309,64'h53c76871dff702a1,64'he1109771607742d1,64'h7456a44b5ed13a7b,
64'h4c594d457ad44a1a,64'h7d9e273027763747,64'hb621e76cc2092f0b,64'h0001fffffffffffe,
64'h07ff0fccdbcb86f9,64'h8649a1cb07daee87,64'hbf45463d8ae17973,64'h2a1021ac5e98bdc2,
64'hfe1caa2492425795,64'h912b7e3e532ae35f,64'had74e568be597f1d,64'hbcdf45f9f477dc17,
64'h3363eb649c7774a6,64'h98ab1f7e5ee24a66,64'hcece8db3789838c8,64'h15650a3d4010f99f,
64'h53beed1873bbfc8c,64'h92b9b98acd77580b,64'hdf66ff35b1ff1777,64'hdf82e404d62e30fd,
64'hfa6d8f66751c4adb,64'h87dc788a902d3360,64'h552731cdaf01e43c,64'h671fbb66d8f2ad83,
64'h6d1fd073c6608d56,64'h8be47576f9b21628,64'h613d0239dbe1be0e,64'h44309b82a25eb5d9,
64'h0230f4a6d2b36bbe,64'h099dc48241d16911,64'h0a029089500d9c6e,64'h0acea559bb2b208b,
64'h1d05d8387169f3a5,64'h8b2464474a3e4e00,64'h376dbe66953f544b,64'hfffff7ff00000801,
64'hfd465cc178e27269,64'h1ec0c3d2a9ebef34,64'h465e9701cdff2977,64'hd86a31ec2a954387,
64'h398e6a0019f8c630,64'hd7fe1019965f1c57,64'he0269bdb2a91de4f,64'hfa557e4125359ca4,
64'h254994d8fda6b29e,64'hc6a5affa1a5d8d82,64'hc7e2c0d4a410a62b,64'ha74851ccd6231195,
64'h466a2184f2d434f3,64'hd7efb2b6890247d9,64'h910c20134791749b,64'h50f69616a595021c,
64'h69b6a05638405835,64'h4436ab982db7e3d1,64'h67c02529367e3b06,64'h16dae05fd5fc6bc5,
64'hd8b3aa69541eac15,64'h752121d084008af8,64'h4f01ddbca741ea4d,64'hb79e92d42fe5a9f3,
64'h192db33abb439844,64'h9e3b4390ffb81506,64'h0884bb9203ba1681,64'ha2b5225df689d3d5,
64'h62ca6a2dd6a250ce,64'hecf139843bb1ba35,64'hb10f3b6b10497853,64'h000ffffffffffff0,
64'h3ff87e66de5c37c8,64'h324d0e5c3ed77434,64'hfa2a31f1570bcb93,64'h50810d63f4c5ee0f,
64'hf0e5512b9212bca1,64'h895bf1f699571af4,64'h6ba72b4af2cbf8e3,64'he6fa2fd4a3bee0b3,
64'h9b1f5b25e3bba52f,64'hc558fbf6f712532c,64'h76746da1c4c1c63a,64'hab2851ea0087ccf8,
64'h9df768c59ddfe45e,64'h95cdcc5a6bbac054,64'hfb37f9b38ff8bbb2,64'hfc17202cb17187e2,
64'hd36c7b3aa8e256d1,64'h3ee3c45881699afc,64'ha9398e6f780f21de,64'h38fddb39c7956c15,
64'h68fe83a133046aad,64'h5f23abbbcd90b13c,64'h09e811d1df0df06d,64'h2184dc1712f5aec6,
64'h1187a536959b5df0,64'h4cee24120e8b4888,64'h5014844a806ce370,64'h56752acdd9590458,
64'he82ec1c38b4f9d28,64'h5923223e51f26ffc,64'hbb6df335a9faa257,64'hffffbfff00004001,
64'hea32e612c7139341,64'hf6061e954f5f79a0,64'h32f4b8106ff94bb6,64'hc3518f6754aa1c32,
64'hcc735001cfc6317f,64'hbff080d2b2f8e2b2,64'h0134dee0548ef271,64'hd2abf21029ace519,
64'h2a4ca6c8ed3594ef,64'h352d7fd6d2ec6c0a,64'h3f1606ab20853152,64'h3a428e6bb1188ca3,
64'h33510c2996a1a796,64'hbf7d95ba48123ec2,64'h8861009e3c8ba4d4,64'h87b4b0b72ca810de,
64'h4db502b4c202c1a5,64'h21b55cc36dbf1e86,64'h3e01294cb3f1d82d,64'hb6d702feafe35e28,
64'hc59d5350a0f560a2,64'ha9090e87200457bd,64'h780eede73a0f5266,64'hbcf496a67f2d4f93,
64'hc96d99d5da1cc220,64'hf1da1c8bfdc0a82c,64'h4425dc901dd0b408,64'h15a912f4b44e9ea3,
64'h16535171b512866d,64'h6789cc28dd8dd1a1,64'h8879db5d824bc293,64'h007fffffffffff80,
64'hffc3f337f2e1be3f,64'h926872e2f6bba19f,64'hd1518f91b85e5c91,64'h84086b21a62f7076,
64'h872a89639095e501,64'h4adf8fb8cab8d79c,64'h5d395a5a965fc715,64'h37d17eac1df70591,
64'hd8fad9331ddd2974,64'h2ac7dfbdb892995a,64'hb3a36d11260e31cd,64'h59428f55043e67bb,
64'hefbb4630eeff22ec,64'hae6e62d75dd6029c,64'hd9bfcda37fc5dd89,64'he0b9016c8b8c3f09,
64'h9b63d9db4712b682,64'hf71e22c50b4cd7df,64'h49cc7380c0790eeb,64'hc7eed9cf3cab60a7,
64'h47f41d0c98235565,64'hf91d5de06c8589de,64'h4f408e8ef86f8368,64'h0c26e0b997ad762f,
64'h8c3d29b4acdaef80,64'h67712092745a443e,64'h80a4225603671b7e,64'hb3a95670cac822be,
64'h41760e235a7ce939,64'hc91911f48f937fde,64'hdb6f99b24fd512b3,64'hfffdffff00020001,
64'h5197309d389c9a01,64'hb030f4b17afbccf9,64'h97a5c0847fca5daf,64'h1a8c7b40a550e18a,
64'h639a80147e318bf2,64'hff84069a97c7158b,64'h09a6f702a4779388,64'h955f90874d6728c2,
64'h5265364869aca777,64'ha96bfeb79763604f,64'hf8b0355a04298a8f,64'hd214735e88c46517,
64'h9a88614db50d3caf,64'hfbecadd74091f60b,64'h430804f5e45d269c,64'h3da585bd654086ec,
64'h6da815a810160d26,64'h0daae61c6df8f42f,64'hf0094a669f8ec167,64'hb6b817fa7f1af13b,
64'h2cea9a8b07ab050a,64'h4848743e0022bde3,64'hc0776f3cd07a932d,64'he7a4b538f96a7c93,
64'h4b6cceb4d0e610fa,64'h8ed0e466ee054159,64'h212ee482ee85a03e,64'had4897a5a274f518,
64'hb29a8b8da8943368,64'h3c4e6149ec6e8d05,64'h43cedaf0125e1494,64'h03fffffffffffc00,
64'hfe1f99c6970df1f1,64'h9343971bb5dd0cf4,64'h8a8c7c93c2f2e482,64'h20435911317b83ac,
64'h39544b2084af2804,64'h56fc7dc855c6bcde,64'he9cad2d6b2fe38a6,64'hbe8bf561efb82c87,
64'hc7d6c99eeee94b9a,64'h563efdeec494cacf,64'h9d1b688e30718e63,64'hca147aaa21f33dd6,
64'h7dda318e77f91759,64'h737316bfeeb014db,64'hcdfe6d21fe2eec42,64'h05c80b6b5c61f841,
64'hdb1ecede3895b40c,64'hb8f1162f5a66bef1,64'h4e639c0803c87756,64'h3f76ce7fe55b0532,
64'h3fa0e866c11aab26,64'hc8eaef0a642c4ee9,64'h7a047479c37c1b3e,64'h613705ccbd6bb178,
64'h61e94da966d77bfc,64'h3b890496a2d221ed,64'h052112b41b38dbec,64'h9d4ab38b564115eb,
64'h0bb0711cd3e749c6,64'h48c88faa7c9bfeea,64'hdb7ccd987ea89592,64'hffefffff00100001,
64'h8cb984ebc4e4d006,64'h8187a590d7de67c3,64'hbd2e0427fe52ed74,64'hd463da052a870c50,
64'h1cd400a6f18c5f8d,64'hfc2034dbbe38ac51,64'h4d37b81523bc9c40,64'haafc843e6b39460c,
64'h9329b2454d653bb6,64'h4b5ff5c1bb1b0273,64'hc581aad7214c5471,64'h90a39afa462328b2,
64'hd4430a71a869e574,64'hdf656ec1048fb051,64'h184027b122e934de,64'hed2c2dec2a04375f,
64'h6d40ad4380b0692d,64'h6d5730e36fc7a178,64'h804a533bfc760b31,64'hb5c0bfd8f8d789d3,
64'h6754d4593d58284f,64'h4243a1f20115ef16,64'h03bb79ec83d49962,64'h3d25a9cecb53e491,
64'h5b6675a8873087ce,64'h7687233b702a0ac4,64'h09772418742d01ef,64'h6a44bd3213a7a8bb,
64'h94d45c7244a19b3b,64'he2730a5063746827,64'h1e76d78292f0a49e,64'h1fffffffffffe000,
64'hf0fcce3bb86f8f81,64'h9a1cb8e1aee8679c,64'h5463e4a21797240c,64'h021ac88a8bdc1d5f,
64'hcaa259052579401f,64'hb7e3ee44ae35e6ee,64'h4e5696bc97f1c529,64'hf45fab147dc16433,
64'h3eb64cfd774a5cca,64'hb1f7ef7824a65676,64'he8db4475838c7314,64'h50a3d5570f99eeaa,
64'heed18c76bfc8bac5,64'h9b98b6027580a6d5,64'h6ff36915f177620a,64'h2e405b5ae30fc208,
64'hd8f676f7c4ada05a,64'hc788b17fd335f783,64'h731ce0421e43baae,64'hfbb674002ad8298f,
64'hfd07433708d5592f,64'h4757785921627742,64'hd023a3d11be0d9ed,64'h09b82e68eb5d8bbd,
64'h0f4a6d4e36bbdfdd,64'hdc4824b616910f67,64'h290895a0d9c6df60,64'hea559c5eb208af54,
64'h5d8388e69f3a4e30,64'h46447d55e4dff74e,64'hdbe66cc9f544ac8a,64'hff7fffff00800001,
64'h65cc27622726802c,64'h0c3d2c8abef33e14,64'he9702144f2976b9b,64'ha31ed02f5438627a,
64'he6a005378c62fc68,64'he101a6e4f1c56281,64'h69bdc0ab1de4e1fe,64'h57e421f859ca305b,
64'h994d922e6b29ddac,64'h5affae0fd8d81396,64'h2c0d56bf0a62a382,64'h851cd7d63119458c,
64'ha2185393434f2b9a,64'hfb2b760e247d8282,64'hc2013d891749a6f0,64'h69616f685021baf1,
64'h6a056a1f05834965,64'h6ab9871e7e3d0bbd,64'h025299e3e3b05984,64'hae05feccc6bc4e93,
64'h3aa6a2cceac14275,64'h121d0f9208af78ae,64'h1ddbcf641ea4cb10,64'he92d4e775a9f2487,
64'hdb33ad4639843e6e,64'hb43919de8150561d,64'h4bb920c3a1680f78,64'h5225e9939d3d45d5,
64'ha6a2e396250cd9d4,64'h1398528a1ba34131,64'hf3b6bc14978524f0,64'h00000000fffeffff,
64'h87e671e4c37c7c01,64'hd0e5c71177433cdc,64'ha31f2512bcb9205e,64'h10d644545ee0eaf8,
64'h5512c82f2bca00f2,64'hbf1f722a71af376b,64'h72b4b5e6bf8e2946,64'ha2fd58aaee0b2191,
64'hf5b267ecba52e64f,64'h8fbf7bc62532b3ab,64'h46da23b31c639899,64'h851eaaba7ccf754e,
64'h768c63bcfe45d621,64'hdcc5b017ac0536a4,64'h7f9b48b28bbb104d,64'h7202dad8187e103f,
64'hc7b3b7c4256d02ca,64'h3c458c0499afbc12,64'h98e70213f21dd56d,64'hddb3a00856c14c71,
64'he83a19bf46aac971,64'h3abbc2cb0b13ba0e,64'h811d1e8edf06cf62,64'h4dc173475aec5de8,
64'h7a536a71b5defee8,64'he24125b6b4887b32,64'h4844ad07ce36faff,64'h52ace2fc90457a99,
64'hec1c4736f9d2717e,64'h3223eab126ffba6e,64'hdf336655aa25644a,64'hfbffffff04000001,
64'h2e613b143934015d,64'h61e96455f799f0a0,64'h4b810a2e94bb5cd1,64'h18f6817fa1c313cb,
64'h350029c36317e339,64'h080d372e8e2b1401,64'h4dee055bef270fed,64'hbf210fc4ce5182d6,
64'hca6c9177594eed5c,64'hd7fd7080c6c09cae,64'h606ab5f953151c0f,64'h28e6beb588ca2c5c,
64'h10c29c9f1a795ccb,64'hd95bb07823ec1409,64'h1009ec4eba4d377a,64'h4b0b7b45810dd785,
64'h502b50fb2c1a4b25,64'h55cc38f6f1e85de5,64'h1294cf1f1d82cc20,64'h702ff66b35e27493,
64'hd5351668560a13a7,64'h90e87c90457bc570,64'heede7b20f5265880,64'h496a73c1d4f92431,
64'hd99d6a37cc21f36a,64'ha1c8cef90a82b0e3,64'h5dc9061f0b407bbe,64'h912f4c9ee9ea2ea6,
64'h35171cb62866ce9b,64'h9cc29450dd1a0988,64'h9db5e0abbc292779,64'h00000007fff7fff8,
64'h3f338f2a1be3e004,64'h872e3891ba19e6da,64'h18f9289ae5c902eb,64'h86b222a2f70757c0,
64'ha896417b5e50078e,64'hf8fb91588d79bb53,64'h95a5af38fc714a2d,64'h17eac55c70590c83,
64'had933f6cd2973271,64'h7dfbde3529959d54,64'h36d11d9ae31cc4c6,64'h28f555d7e67baa6c,
64'hb4631deaf22eb105,64'he62d80c36029b51a,64'hfcda45975dd88265,64'h9016d6c3c3f081f5,
64'h3d9dbe272b68164a,64'he22c6025cd7de08f,64'hc73810a390eeab64,64'hed9d0048b60a6382,
64'h41d0ce0135564b81,64'hd5de1659589dd06f,64'h08e8f47af8367b0c,64'h6e0b9a3cd762ef3e,
64'hd29b5390aef7f73d,64'h12092dbca443d989,64'h4225684071b7d7f6,64'h956717e6822bd4c6,
64'h60e239bece938be9,64'h911f558a37fdd36f,64'hf99b32b3512b224a,64'hdfffffff20000001,
64'h7309d8a2c9a00ae7,64'h0f4b22b2bccf84fd,64'h5c085176a5dae686,64'hc7b40bfd0e189e58,
64'ha8014e1c18bf19c7,64'h4069b9747158a008,64'h6f702ae179387f66,64'hf9087e2b728c16ab,
64'h53648bc0ca776ada,64'hbfeb840c3604e56a,64'h0355afcd98a8e075,64'h4735f5ad465162df,
64'h8614e4f8d3cae658,64'hcadd83c71f60a042,64'h804f6275d269bbd0,64'h585bda2e086ebc26,
64'h815a87db60d25926,64'hae61c7b98f42ef26,64'h94a678f8ec166100,64'h817fb35caf13a495,
64'ha9a8b348b0509d32,64'h8743e4862bde2b7c,64'h76f3d90ea932c3f9,64'h4b539e10a7c92186,
64'hcceb51c4610f9b4a,64'h0e4677cd54158713,64'hee4830fa5a03ddee,64'h897a64fb4f51752c,
64'ha8b8e5b2433674d7,64'he614a28ae8d04c3c,64'hedaf0561e1493bc4,64'h0000003fffbfffc0,
64'hf99c7951df1f001f,64'h3971c491d0cf36cc,64'hc7c944d72e481758,64'h3591151bb83abdfc,
64'h44b20bdff2803c6b,64'hc7dc8acb6bcdda91,64'had2d79cbe38a5164,64'hbf562ae382c86418,
64'h6c99fb6b94b99383,64'hefdef1ac4cacea9d,64'hb688ecd818e6262f,64'h47aaaec033dd535f,
64'ha318ef5c91758823,64'h316c0622014da8c9,64'he6d22cc1eec41321,64'h80b6b6221f840fa4,
64'hecedf13a5b40b24f,64'h116301356bef0471,64'h39c0852287755b1a,64'h6ce8024cb0531c09,
64'h0e86700baab25c06,64'haef0b2d0c4ee8372,64'h4747a3d7c1b3d860,64'h705cd1e9bb1779ed,
64'h94da9c8b77bfb9e2,64'h90496de5221ecc48,64'h112b42058dbebfae,64'hab38bf38115ea62c,
64'h0711cdf9749c5f45,64'h88faac55bfee9b74,64'hccd995a189591249,64'h0000000000000001
};
  //------------------------
  // 1024
  //------------------------
  localparam [2*1024-1:0][63:0] NTT_GF64_BWD_N1024_PHI_L = {
64'h7a591595e67c27e8,64'h3da05fee70c4f2ba,64'h034dcba58ac5003e,64'hc843f1629460b551,
64'hff5c2066b0272b4b,64'h39afad6c328b16f6,64'h56ec1e3efb05020a,64'hc2ded1724375e12e,
64'h730e3dd17a17792b,64'h0bfd9ae9789d24a4,64'h3a1f24355ef15bdc,64'h5a9cf0873e490c2e,
64'h7233be6aa0ac3898,64'h4bd327de7a8ba95c,64'h30a5145e468261d9,64'h000001fffdfffe00,
64'hcb8e248f8679b65f,64'hac88a8dec1d5efdf,64'h3ee456615e6ed482,64'hfab15721164320bb,
64'h7ef78d69656754e1,64'h3d5576039eea9af6,64'h8b6031110a6d4647,64'h05b5b114fc207d1c,
64'h8b1809ab5f782388,64'h674012688298e045,64'h7785968b27741b8b,64'h82e68f50d8bbcf65,
64'h824b6f2d10f6623c,64'h59c5f9c58af5315b,64'h47d562b1ff74db9c,64'h0000000000000008,
64'hd2c8acb233e13f3d,64'hed02ff74862795cf,64'h1a6e5d2c562801f0,64'h421f8b1aa305aa82,
64'hfae1033c81395a51,64'hcd7d6b629458b7af,64'hb760f1f9d828104e,64'h16f68b981baf096a,
64'h9871ee8ed0bbc955,64'h5fecd74bc4e92520,64'hd0f921abf78adedf,64'hd4e7843bf248616e,
64'h919df3580561c4bd,64'h5e993ef5d45d4ade,64'h8528a2f334130ec7,64'h00000fffeffff000,
64'h5c71248233cdb2f2,64'h644546fb0eaf7ef3,64'hf722b30bf376a40f,64'hd58ab90fb21905d1,
64'hf7bc6b4e2b3aa705,64'heaabb01df754d7af,64'h5b01888c536a3234,64'h2dad88a7e103e8e0,
64'h58c04d5efbc11c3c,64'h3a00934714c70225,64'hbc2cb45c3ba0dc55,64'h17347a8ac5de7b24,
64'h125b796c87b311dc,64'hce2fce2e57a98ad6,64'h3eab1591fba6dcde,64'h0000000000000040,
64'h964565979f09f9e2,64'h6817fbab313cae71,64'hd372e962b1400f80,64'h10fc58d7182d540e,
64'hd70819eb09cad281,64'h6beb5b1aa2c5bd72,64'hbb078fd3c140826b,64'hb7b45cc0dd784b50,
64'hc38f747a85de4aa4,64'hff66ba60274928fe,64'h87c90d65bc56f6f2,64'ha73c21e592430b6a,
64'h8cef9ac42b0e25e4,64'hf4c9f7b0a2ea56ee,64'h2945179da0987634,64'h00007fff7fff8000,
64'he38924139e6d978e,64'h222a37db757bf795,64'hb91598669bb52071,64'hac55c88390c82e82,
64'hbde35a7859d53821,64'h555d80f6baa6bd71,64'hd80c44649b51919e,64'h6d6c4540081f46ff,
64'hc6026af9de08e1de,64'hd0049a39a6381127,64'he165a2e6dd06e2a3,64'hb9a3d4562ef3d920,
64'h92dbcb643d988ee0,64'h717e7178bd4c56aa,64'hf558ac90dd36e6ef,64'h0000000000000200,
64'hb22b2cc0f84fcf0c,64'h40bfdd5c89e57385,64'h9b974b1b8a007bfa,64'h87e2c6b8c16aa070,
64'hb840cf5e4e569402,64'h5f5ad8d8162deb8d,64'hd83c7ea30a041353,64'hbda2e60bebc25a7b,
64'h1c7ba3da2ef2551a,64'hfb35d3083a4947e9,64'h3e486b31e2b7b78c,64'h39e10f3192185b4b,
64'h677cd62558712f1c,64'ha64fbd8c1752b769,64'h4a28bcee04c3b19f,64'h0003fffbfffc0000,
64'h1c4920a3f36cbc69,64'h1151bedcabdfbca7,64'hc8acc339dda90383,64'h62ae44218641740b,
64'hef1ad3c7cea9c103,64'haaec07b7d535eb86,64'hc062232ada8c8cea,64'h6b622a0340fa37f5,
64'h301357d4f0470eea,64'h8024d1d331c08932,64'h0b2d173de8371511,64'hcd1ea2b6779ec8fb,
64'h96de5b25ecc476fc,64'h8bf38bc8ea62b54d,64'haac5648de9b73771,64'h0000000000001000,
64'h9159660cc27e785b,64'h05feeae64f2b9c26,64'hdcba58e05003dfcc,64'h3f1635ca0b55037c,
64'hc2067af772b4a00b,64'hfad6c6c2b16f5c66,64'hc1e3f51e50209a92,64'hed1730645e12d3d3,
64'he3dd1ed17792a8d0,64'hd9ae9848d24a3f41,64'hf243599015bdbc5f,64'hcf08798d90c2da57,
64'h3be6b12dc38978dd,64'h327dec65ba95bb43,64'h5145e772261d8cf6,64'h001fffdfffe00000,
64'he249051f9b65e348,64'h8a8df6e55efde538,64'h456619d4ed481c12,64'h1572210f320ba055,
64'h78d69e45754e0811,64'h57603dc3a9af5c2b,64'h0311195cd464674a,64'h5b11501d07d1bfa5,
64'h809abea88238774f,64'h01268e9d8e04498c,64'h5968b9ef41b8a888,64'h68f515b9bcf647d2,
64'hb6f2d9336623b7dc,64'h5f9c5e4b5315aa64,64'h562b24744db9bb83,64'h0000000000008000,
64'h8acb306a13f3c2d4,64'h2ff75732795ce130,64'he5d2c708801efe5a,64'hf8b1ae515aa81bdf,
64'h1033d7c195a50052,64'hd6b6361c8b7ae329,64'h0f1fa8f88104d48a,64'h68b98329f0969e91,
64'h1ee8f692bc954679,64'hcd74c24c9251fa02,64'h921acc87adede2f1,64'h7843cc728616d2b2,
64'hdf35896f1c4bc6e7,64'h93ef632ed4adda17,64'h8a2f3b9330ec67ae,64'h00fffeffff000000,
64'h12482903db2f1a39,64'h546fb72ef7ef29bc,64'h2b30cea96a40e08e,64'hab910879905d02a8,
64'hc6b4f22eaa704085,64'hbb01ee1f4d7ae156,64'h1888cae6a3233a50,64'hd88a80ea3e8dfd26,
64'h04d5f54811c3ba74,64'h093474ec70224c60,64'hcb45cf7c0dc5443e,64'h47a8add0e7b23e8d,
64'hb796c9a0311dbedb,64'hfce2f25c98ad531e,64'hb15923a46dcddc16,64'h0000000000040000,
64'h565983549f9e169c,64'h7fbab994cae7097f,64'h2e96384b00f7f2c9,64'hc58d7291d540def1,
64'h819ebe0cad280290,64'hb5b1b0ea5bd71942,64'h78fd47c40826a450,64'h45cc195284b4f485,
64'hf747b495e4aa33c8,64'h6ba6126a928fd00a,64'h90d664416f6f1784,64'hc21e639730b6958d,
64'hf9ac4b7ee25e3732,64'h9f7b197aa56ed0b4,64'h5179dc9d87633d6c,64'h07fff7fff8000000,
64'h9241481ed978d1c8,64'ha37db979bf794dde,64'h5986754c5207046f,64'h5c8843d182e8153b,
64'h35a7917b53820422,64'hd80f70ff6bd70aab,64'hc44657351919d280,64'hc4540757f46fe92a,
64'h26afaa408e1dd3a0,64'h49a3a76381126300,64'h5a2e7be66e2a21ea,64'h3d456e893d91f466,
64'hbcb64d0688edf6d3,64'he71792ebc56a98e9,64'h8ac91d286e6ee0ab,64'h0000000000200000,
64'hb2cc1aa6fcf0b4de,64'hfdd5cca957384bf5,64'h74b1c25907bf9647,64'h2c6b9494aa06f782,
64'h0cf5f0696940147c,64'had8d8757deb8ca0b,64'hc7ea3e234135227d,64'h2e60ca9625a7a426,
64'hba3da4b625519e39,64'h5d309357947e804d,64'h86b3220f7b78bc1c,64'h10f31cbf85b4ac62,
64'hcd625bfe12f1b989,64'hfbd8cbd92b76859c,64'h8bcee4ee3b19eb5e,64'h3fffbfffc0000000,
64'h920a40facbc68e3c,64'h1bedcbd2fbca6eeb,64'hcc33aa6490382376,64'he4421e8e1740a9d6,
64'had3c8bdb9c10210f,64'hc07b88015eb85552,64'h2232b9aec8ce93fa,64'h22a03ac5a37f494a,
64'h357d520570ee9cff,64'h4d1d3b1e089317fe,64'hd173df3571510f4e,64'hea2b744aec8fa32f,
64'he5b26839476fb693,64'h38bc97652b54c741,64'h5648e94773770554,64'h0000000001000000,
64'h9660d53ce785a6eb,64'heeae6551b9c25fa1,64'ha58e12cb3dfcb235,64'h635ca4a65037bc0f,
64'h67af834b4a00a3e0,64'h6c6c3ac3f5c65053,64'h3f51f12009a913e2,64'h730654b22d3d212f,
64'hd1ed25b62a8cf1c3,64'he9849abea3f40266,64'h3599107fdbc5e0dc,64'h8798e5fc2da56310,
64'h6b12dff6978dcc42,64'hdec65ed05bb42cd9,64'h5e772775d8cf5aec,64'hfffdfffeffffffff,
64'h905207da5e3471dc,64'hdf6e5e97de537758,64'h619d532a81c11baa,64'h2210f477ba054ea9,
64'h69e45ee1e0810873,64'h03dc4010f5c2aa8a,64'h1195cd7746749fcf,64'h1501d62e1bfa4a4f,
64'habea902c8774e7f7,64'h68e9d8f24498bfee,64'h8b9ef9b18a887a6a,64'h515ba25e647d1971,
64'h2d9341d13b7db491,64'hc5e4bb2a5aa63a07,64'hb2474a3d9bb82a9e,64'h0000000008000000,
64'hb306a9eb3c2d3754,64'h75732a94ce12fd01,64'h2c70965eefe591a3,64'h1ae5253581bde075,
64'h3d7c1a5d50051efd,64'h6361d622ae328295,64'hfa8f89014d489f0f,64'h9832a59469e90975,
64'h8f692db754678e12,64'h4c24d5fc1fa01329,64'hacc883ffde2f06df,64'h3cc72fe56d2b187c,
64'h5896ffb7bc6e620d,64'hf632f688dda166c2,64'hf3b93bb0c67ad75e,64'hffeffffefffffff1,
64'h82903ed6f1a38edc,64'hfb72f4c4f29bbaba,64'h0cea99570e08dd4d,64'h1087a3bed02a7547,
64'h4f22f71204084395,64'h1ee20087ae155450,64'h8cae6bba33a4fe78,64'ha80eb170dfd25278,
64'h5f5481693ba73fb3,64'h474ec79524c5ff6d,64'h5cf7cd905443d34c,64'h8add12f523e8cb86,
64'h6c9a0e8adbeda487,64'h2f25d958d531d032,64'h923a51f1ddc154eb,64'h0000000040000000,
64'h98354f5ee169ba9b,64'hab9954a97097e805,64'h6384b2f87f2c8d17,64'hd72929ac0def03a8,
64'hebe0d2eb8028f7e7,64'h1b0eb118719414a5,64'hd47c48116a44f871,64'hc1952ca74f484ba4,
64'h7b496dbea33c708c,64'h6126afe2fd009946,64'h66442003f17836f3,64'he6397f2c6958c3df,
64'hc4b7fdbfe3731066,64'hb197b44ded0b3609,64'h9dc9dd8d33d6bae9,64'hff7ffffeffffff81,
64'h1481f6bb8d1c76dc,64'hdb97a62e94ddd5c9,64'h6754cab87046ea68,64'h843d1df68153aa38,
64'h7917b89220421ca6,64'hf710043d70aaa280,64'h65735dd59d27f3bc,64'h40758b8bfe9293bb,
64'hfaa40b4bdd39fd96,64'h3a763cab262ffb66,64'he7be6c84a21e9a5e,64'h56e897ad1f465c2c,
64'h64d07459df6d2435,64'h792ecac7a98e818f,64'h91d28f92ee0aa754,64'h0000000200000000,
64'hc1aa7afb0b4dd4d4,64'h5ccaa55084bf4023,64'h1c2597c6f96468b5,64'hb9494d666f781d3a,
64'h5f0697630147bf31,64'hd87588c38ca0a528,64'ha3e240915227c382,64'h0ca965407a425d1a,
64'hda4b6df819e3845d,64'h09357f1ae804ca2d,64'h322100228bc1b795,64'h31cbf96a4ac61ef1,
64'h25bfee051b98832a,64'h8cbda2746859b043,64'hee4eec6d9eb5d744,64'hfbfffffefffffc01,
64'ha40fb5dc68e3b6e0,64'hdcbd317aa6eeae42,64'h3aa655c68237533d,64'h21e8efb80a9d51bc,
64'hc8bdc4940210e52d,64'hb88021f2855513f9,64'h2b9aeeafe93f9ddd,64'h03ac5c61f4949dd6,
64'hd5205a65e9cfeca9,64'hd3b1e55a317fdb2f,64'h3df3642c10f4d2e9,64'hb744bd6afa32e15e,
64'h2683a2d1fb6921a5,64'hc97656404c740c75,64'h8e947c9b70553a9c,64'h0000001000000000,
64'h0d53d7de5a6ea69a,64'he6552a8625fa0116,64'he12cbe37cb2345a8,64'hca4a6b387bc0e9cb,
64'hf834bb1a0a3df986,64'hc3ac46226505293a,64'h1f12048f913e1c0b,64'h654b2a03d212e8d0,
64'hd25b6fc6cf1c22e2,64'h49abf8d740265168,64'h910801155e0dbca7,64'h8e5fcb535630f787,
64'h2dff7029dcc4194f,64'h65ed13a742cd8214,64'h72776373f5aeba19,64'hdffffffeffffe001,
64'h207daee8471db6fb,64'he5e98bdb3775720a,64'hd532ae3511ba99e7,64'h0f477dc154ea8ddf,
64'h45ee24a610872962,64'hc4010f992aa89fc3,64'h5cd7758049fceee7,64'h1d62e30fa4a4eeb0,
64'ha902d3354e7f6542,64'h9d8f2ad78bfed972,64'hef9b216187a69747,64'hba25eb5cd1970aeb,
64'h341d1690db490d27,64'h4bb2b20863a063a2,64'h74a3e4df82a9d4dc,64'h0000008000000000,
64'h6a9ebef2d37534d0,64'h32a954382fd008a9,64'h0965f1c5591a2d39,64'h525359c9de074e52,
64'hc1a5d8d751efcc29,64'h1d623119282949ca,64'hf890247c89f0e058,64'h2a5950219097467d,
64'h92db7e3c78e1170a,64'h4d5fc6bc01328b3e,64'h884008aef06de534,64'h72fe5a9eb187bc34,
64'h6ffb814fe620ca77,64'h2f689d3d166c109d,64'h93bb1ba2ad75d0c5,64'hfffffffdffff0002,
64'h03ed774338edb7d7,64'h2f4c5ee0bbab9049,64'ha99571ae8dd4cf32,64'h7a3bee0aa7546ef8,
64'h2f71253284394b0e,64'h20087ccf5544fe12,64'he6bbac044fe77736,64'heb17187d25277580,
64'h481699af73fb2a0b,64'hec7956c05ff6cb8c,64'h7cd90b133d34ba31,64'hd12f5aeb8cb85753,
64'ha0e8b487da486937,64'h5d9590451d031d0e,64'ha51f26ff154ea6dd,64'h0000040000000000,
64'h54f5f7999ba9a67d,64'h954aa1c27e804547,64'h4b2f8e2ac8d169c8,64'h929ace50f03a728e,
64'h0d2ec6c08f7e6142,64'heb1188c9414a4e50,64'hc48123eb4f8702b9,64'h52ca810d84ba33e7,
64'h96dbf1e7c708b84c,64'h6afe35e2099459ee,64'h4200457b836f299c,64'h97f2d4f88c3de19d,
64'h7fdc0a82310653b5,64'h7b44e9e9b36084e7,64'h9dd8dd196bae8624,64'hfffffff6fff80009,
64'h1f6bba19c76dbeb8,64'h7a62f706dd5c8247,64'h4cab8d796ea6798b,64'hd1df70583aa377bd,
64'h7b89299521ca586f,64'h0043e67baa27f08f,64'h35dd60297f3bb9a9,64'h58b8c3f0293babf9,
64'h40b4cd7d9fd95056,64'h63cab609ffb65c59,64'he6c8589ce9a5d185,64'h897ad76265c2ba92,
64'h0745a443d24349b3,64'hecac822ae818e86e,64'h28f937fdaa7536e3,64'h0000200000000000,
64'ha7afbccedd4d33e6,64'haa550e17f4022a34,64'h597c7158468b4e3e,64'h94d6728b81d3946c,
64'h697636047bf30a10,64'h588c46510a527279,64'h24091f607c3815c2,64'h9654086e25d19f36,
64'hb6df8f423845c25c,64'h57f1af134ca2cf6d,64'h10022bde1b794cde,64'hbf96a7c861ef0ce4,
64'hfee0541488329da5,64'hda274f509b042735,64'heec6e8cf5d74311c,64'hffffffbeffc00041,
64'hfb5dd0ce3b6df5c0,64'hd317b839eae41235,64'h655c6bcd7533cc56,64'h8efb82c7d51bbde2,
64'hdc494cac0e52c375,64'h021f33dd513f8478,64'haeeb014cf9ddcd47,64'hc5c61f8349dd5fc6,
64'h05a66beefeca82ae,64'h1e55b052fdb2e2c5,64'h3642c4ee4d2e8c21,64'h4bd6bb172e15d48c,
64'h3a2d221e921a4d98,64'h6564115e40c74369,64'h47c9bfee53a9b717,64'h0001000000000000,
64'h3d7de67bea699f2b,64'h52a870c4a011519b,64'hcbe38ac4345a71ee,64'ha6b394600e9ca35c,
64'h4bb1b026df98507d,64'hc462328a529393c6,64'h2048fb04e1c0ae0f,64'hb2a043752e8cf9ac,
64'hb6fc7a16c22e12db,64'hbf8d789c65167b66,64'h80115ef0dbca66f0,64'hfcb53e480f78671b,
64'hf702a0ab4194ed21,64'hd13a7a8ad82139a2,64'h76374681eba188d9,64'hfffffdfefe000201,
64'hdaee8678db6fadf9,64'h98bdc1d5572091a2,64'h2ae35e6ea99e62ad,64'h77dc1642a8ddef0c,
64'he24a656672961ba2,64'h10f99eea89fc23c0,64'h77580a6cceee6a33,64'h2e30fc204eeafe2a,
64'h2d335f77f6541570,64'hf2ad8297ed971628,64'hb216277369746107,64'h5eb5d8bb70aea45e,
64'hd16910f590d26cbf,64'h2b208af5063a1b45,64'h3e4dff749d4db8b6,64'h0008000000000000,
64'hebef33e0534cf957,64'h95438627008a8cd6,64'h5f1c5627a2d38f6a,64'h359ca30574e51adb,
64'h5d8d8138fcc283e6,64'h23119458949c9e2a,64'h0247d8280e057077,64'h95021bae7467cd5b,
64'hb7e3d0bb117096d3,64'hfc6bc4e828b3db2b,64'h008af78ade53377c,64'he5a9f2477bc338d1,
64'hb81505610ca76901,64'h89d3d45cc109cd0a,64'hb1ba34125d0c46c5,64'hffffeffef0001001,
64'hd77433ccdb7d6fc2,64'hc5ee0eaeb9048d0c,64'h571af3764cf31567,64'hbee0b21846ef785d,
64'h12532b3a94b0dd09,64'h87ccf7544fe11e00,64'hbac0536977735195,64'h7187e1037757f14f,
64'h699afbc0b2a0ab7f,64'h956c14c66cb8b139,64'h90b13ba04ba30833,64'hf5aec5dd857522ee,
64'h8b4887b2869365f2,64'h590457a931d0da27,64'hf26ffba5ea6dc5af,64'h0040000000000000,
64'h5f799f099a67cab1,64'haa1c313c045466ac,64'hf8e2b13f169c7b4e,64'hace5182ca728d6d7,
64'hec6c09c9e6141f2e,64'h188ca2c5a4e4f14f,64'h123ec140702b83b8,64'ha810dd77a33e6ad4,
64'hbf1e85dd8b84b693,64'he35e2748459ed951,64'h0457bc56f299bbe0,64'h2d4f9242de19c681,
64'hc0a82b0d653b4803,64'h4e9ea2ea084e684c,64'h8dd1a097e8623623,64'hffff7ffe80008001,
64'hbba19e6cdbeb7e0a,64'h2f70757bc824685a,64'hb8d79bb46798ab36,64'hf70590c7377bc2e3,
64'h929959d4a586e848,64'h3e67baa67f08effc,64'hd6029b50bb9a8ca3,64'h8c3f081ebabf8a75,
64'h4cd7de0895055bf5,64'hab60a63765c589c4,64'h8589dd065d184194,64'had762ef32ba91769,
64'h5a443d98349b2f8c,64'hc822bd4b8e86d136,64'h937fdd36536e2d71,64'h0200000000000000,
64'hfbccf84ed33e5586,64'h50e189e522a3355b,64'hc71589ffb4e3da69,64'h6728c16a3946b6b3,
64'h63604e5630a0f969,64'hc465162d27278a78,64'h91f60a03815c1dc0,64'h4086ebc219f3569b,
64'hf8f42ef15c25b493,64'h1af13a492cf6ca81,64'h22bde2b794cddf00,64'h6a7c9217f0ce3407,
64'h0541587129da4012,64'h74f517524273425e,64'h6e8d04c34311b114,64'hfffbfffb00040001,
64'hdd0cf36bdf5bf04b,64'h7b83abdf412342cf,64'hc6bcdda83cc559ab,64'hb82c8640bbde1711,
64'h94cacea92c37423c,64'hf33dd534f8477fdf,64'hb014da8bdcd46512,64'h61f840f9d5fc53a4,
64'h66bef046a82adfa6,64'h5b0531c02e2c4e1b,64'h2c4ee836e8c20c9c,64'h6bb1779e5d48bb43,
64'hd221ecc3a4d97c5e,64'h4115ea62743689aa,64'h9bfee9b69b716b84,64'h1000000000000000,
64'hde67c27d99f2ac29,64'h870c4f2b1519aad6,64'h38ac5003a71ed342,64'h39460b54ca35b595,
64'h1b0272b48507cb45,64'h2328b16f393c53ba,64'h8fb050200ae0edfc,64'h04375e12cf9ab4d6,
64'hc7a17791e12da491,64'hd789d24967b65408,64'h15ef15bda66ef7ff,64'h53e490c28671a035,
64'h2a0ac3894ed20090,64'ha7a8ba95139a12ed,64'h7468261d188d889d,64'hffdfffdf00200001,
64'he8679b64fadf8252,64'hdc1d5efd091a1675,64'h35e6ed47e62acd52,64'hc164320adef0b883,
64'ha656754d61ba11dc,64'h99eea9aec23bfef1,64'h80a6d463e6a3288b,64'h0fc207d1afe29d1d,
64'h35f782384156fd2d,64'hd8298e03716270d6,64'h627741b8461064df,64'h5d8bbcf5ea45da15,
64'h910f662326cbe2ea,64'h08af5315a1b44d4e,64'hdff74db8db8b5c1c,64'h8000000000000000,
64'hf33e13f2cf956142,64'h3862795ca8cd56ac,64'hc562801e38f69a0f,64'hca305aa751adaca7,
64'hd81395a4283e5a28,64'h19458b7ac9e29dcf,64'h7d82810457076fdc,64'h21baf0967cd5a6b0,
64'h3d0bbc95096d2482,64'hbc4e92513db2a03a,64'haf78aded3377bff8,64'h9f248616338d01a6,
64'h50561c4b7690047f,64'h3d45d4ad9cd09763,64'ha34130ebc46c44e5,64'hfefffeff01000001,
64'h433cdb2ed6fc1289,64'he0eaf7ee48d0b3a2,64'haf376a4031566a8f,64'h0b21905cf785c412,
64'h32b3aa700dd08edb,64'hcf754d7a11dff784,64'h0536a32335194454,64'h7e103e8d7f14e8e8,
64'hafbc11c30ab7e967,64'hc14c70218b1386aa,64'h13ba0dc5308326f5,64'hec5de7b1522ed0a6,
64'h887b311d365f174c,64'h457a98ad0da26a70,64'hffba6dccdc5ae0da,64'h00000003fffffffc,
64'h99f09f9d7cab0a09,64'hc313cae6466ab55f,64'h2b1400f7c7b4d072,64'h5182d5408d6d6532,
64'hc09cad2741f2d13a,64'hca2c5bd64f14ee78,64'hec140825b83b7edd,64'h0dd784b4e6ad357f,
64'he85de4a94b69240f,64'he274928eed9501cb,64'h7bc56f6e9bbdffbb,64'hf92430b59c680d2c,
64'h82b0e25db48023f6,64'hea2ea56de684bb17,64'h1a09876323622723,64'hf7fff7ff08000001,
64'h19e6d978b7e09446,64'h0757bf7946859d09,64'h79bb52068ab35473,64'h590c82e7bc2e2090,
64'h959d53816e8476d7,64'h7baa6bd68effbc1a,64'h29b51919a8ca22a0,64'hf081f46ef8a7473d,
64'h7de08e1d55bf4b33,64'h0a638112589c354a,64'h9dd06e29841937a8,64'h62ef3d9191768529,
64'h43d988edb2f8ba5c,64'h2bd4c56a6d13537e,64'hfdd36e6de2d706c9,64'h0000001fffffffe0,
64'hcf84fcefe5585044,64'h189e57383355aaf2,64'h58a007bf3da6838f,64'h8c16aa066b6b298e,
64'h04e569400f9689ca,64'h5162deb878a773ba,64'h60a04134c1dbf6e1,64'h6ebc25a73569abf8,
64'h42ef25515b492071,64'h13a4947e6ca80e51,64'hde2b7b77ddeffdd5,64'hc92185b3e3406959,
64'h158712f1a4011fac,64'h51752b763425d8b1,64'hd04c3b191b113918,64'hbfffbfff40000001,
64'hcf36cbc5bf04a230,64'h3abdfbca342ce848,64'hcdda9037559aa395,64'hc864173fe171047e,
64'hacea9c0f7423b6b4,64'hdd535eb777fde0cd,64'h4da8c8ce465114ff,64'h840fa37ec53a39e1,
64'hef0470edadfa5995,64'h531c0892c4e1aa50,64'hee83715020c9bd3c,64'h1779ec8f8bb42945,
64'h1ecc476f97c5d2de,64'h5ea62b54689a9bef,64'hee9b737616b83641,64'h000000ffffffff00,
64'h7c27e7852ac2821a,64'hc4f2b9c19aad5790,64'hc5003dfbed341c76,64'h60b550375b594c6c,
64'h272b4a007cb44e50,64'h8b16f5c5c53b9dce,64'h050209a90edfb705,64'h75e12d3cab4d5fbd,
64'h17792a8cda490386,64'h9d24a3f365407288,64'hf15bdbc4ef7feea2,64'h490c2da51a034ac2,
64'hac38978d2008fd60,64'h8ba95bb3a12ec586,64'h8261d8ced889c8ba,64'hfffdffff00000003,
64'h79b65e33f825117a,64'hd5efde52a167423f,64'h6ed481c0acd51ca2,64'h4320ba050b8823ea,
64'h6754e080a11db59b,64'hea9af5c1bfef0662,64'h6d4646743288a7f6,64'h207d1bfa29d1cf04,
64'h782387746fd2cca1,64'h98e04498270d527e,64'h741b8a88064de9d9,64'hbbcf647c5da14a28,
64'hf6623b7cbe2e96f0,64'hf5315aa544d4df76,64'h74db9bb7b5c1b201,64'h000007fffffff800,
64'he13f3c2c561410cd,64'h2795ce12d56abc7a,64'h2801efe569a0e3aa,64'h05aa81bddaca635d,
64'h395a5004e5a2727f,64'h58b7ae3229dcee6c,64'h28104d4876fdb828,64'haf0969e85a6afde5,
64'hbbc95466d2481c30,64'he9251f9f2a03943c,64'h8adede2e7bff7509,64'h48616d2ad01a560e,
64'h61c4bc6e0047eafb,64'h5d4adda109762c2c,64'h130ec67ac44e45cc,64'hffefffff00000011,
64'hcdb2f1a2c1288bcd,64'haf7ef29b0b3a11f2,64'h76a40e0866a8e50d,64'h1905d02a5c411f4e,
64'h3aa7040808edacd5,64'h54d7ae14ff783309,64'h6a3233a494453fad,64'h03e8dfd24e8e781f,
64'hc11c3ba67e966505,64'hc70224c5386a93ec,64'ha0dc5443326f4ec5,64'hde7b23e7ed0a513b,
64'hb311dbecf174b779,64'ha98ad53126a6fba9,64'ha6dcddc0ae0d9005,64'h00003fffffffc000,
64'h09f9e169b0a08661,64'h3cae7097ab55e3cf,64'h400f7f2c4d071d4f,64'h2d540deed6531ae8,
64'hcad280282d1393f7,64'hc5bd71934ee7735e,64'h40826a44b7edc13f,64'h784b4f47d357ef23,
64'hde4aa33b9240e17b,64'h4928fd00501ca1d9,64'h56f6f177dffba844,64'h430b695880d2b06e,
64'h0e25e373023f57d5,64'hea56ed0a4bb1615e,64'h987633d622722e60,64'hff7fffff00000081,
64'h6d978d1c09445e62,64'h7bf794dd59d08f8b,64'hb520704635472865,64'hc82e8152e208fa70,
64'hd5382041476d66a7,64'ha6bd70a9fbc19846,64'h51919d27a229fd65,64'h1f46fe927473c0f8,
64'h08e1dd39f4b32822,64'h3811262fc3549f5a,64'h06e2a21e937a7623,64'hf3d91f45685289d2,
64'h988edf6c8ba5bbc3,64'h4c56a98e3537dd43,64'h36e6ee0a706c8023,64'h0001fffffffe0000,
64'h4fcf0b4d85043308,64'he57384be5aaf1e77,64'h007bf9646838ea76,64'h6aa06f77b298d73f,
64'h56940147689c9fb2,64'h2deb8ca0773b9aea,64'h04135227bf6e09f6,64'hc25a7a419abf7915,
64'hf25519e292070bd2,64'h4947e80480e50ec6,64'hb7b78bc0ffdd421e,64'h185b4ac60695836e,
64'h712f1b9811fabea8,64'h52b768595d8b0ae9,64'hc3b19eb5139172fc,64'hfbffffff00000401,
64'h6cbc68e34a22f30d,64'hdfbca6edce847c55,64'ha9038236aa394323,64'h41740a9d1047d37a,
64'ha9c102103b6b3532,64'h35eb8554de0cc22b,64'h8c8ce93f114feb26,64'hfa37f493a39e07c0,
64'h470ee9cfa5994110,64'hc089317f1aa4facf,64'h371510f49bd3b118,64'h9ec8fa3242944e89,
64'hc476fb685d2dde14,64'h62b54c73a9beea16,64'hb737705483640117,64'h000ffffffff00000,
64'h7e785a6e2821983e,64'h2b9c25f9d578f3b1,64'h03dfcb2341c753b0,64'h55037bc094c6b9f5,
64'hb4a00a3d44e4fd8e,64'h6f5c6504b9dcd74f,64'h209a913dfb704fb0,64'h12d3d212d5fbc8a2,
64'h92a8cf1b90385e89,64'h4a3f40260728762e,64'hbdbc5e0cfeea10eb,64'hc2da563034ac1b70,
64'h8978dcc38fd5f53d,64'h95bb42ccec585746,64'h1d8cf5ae9c8b97da,64'hdfffffff00002001,
64'h65e3471d51179865,64'hfde537747423e2a2,64'h481c11ba51ca1913,64'h0ba054ea823e9bce,
64'h4e081086db59a98b,64'haf5c2aa7f0661157,64'h646749fc8a7f592c,64'hd1bfa4a41cf03df9,
64'h38774e7f2cca087e,64'h04498bfed527d672,64'hb8a887a5de9d88bf,64'hf647d19614a27444,
64'h23b7db48e96ef09a,64'h15aa63a04df750ad,64'hb9bb82a91b2008b3,64'h007fffffff800000,
64'hf3c2d374410cc1ed,64'h5ce12fcfabc79d87,64'h1efe591a0e3a9d80,64'ha81bde06a635cfa6,
64'ha50051ef2727ec6b,64'h7ae32828cee6ba75,64'h04d489f0db827d7f,64'h969e9096afde4510,
64'h954678e081c2f444,64'h51fa01323943b16e,64'hede2f06cf7508753,64'h16d2b187a560db7a,
64'h4bc6e6207eafa9e4,64'hadda166b62c2ba2c,64'hec67ad74e45cbed0,64'hfffffffe00010002,
64'h2f1a38ed88bcc325,64'hef29bbaaa11f1509,64'h40e08dd48e50c896,64'h5d02a75411f4de70,
64'h70408438dacd4c56,64'h7ae1554483308ab3,64'h233a4fe753fac95d,64'h8dfd2526e781efc2,
64'hc3ba73fa665043ef,64'h224c5ff6a93eb390,64'hc5443d33f4ec45f3,64'hb23e8cb7a513a219,
64'h1dbeda484b7784cf,64'had531d026fba8568,64'hcddc154dd9004593,64'h03fffffffc000000,
64'h9e169ba908660f61,64'he7097e7f5e3cec36,64'hf7f2c8d071d4ec00,64'h40def03a31ae7d2b,
64'h28028f7e393f6353,64'hd71941497735d3a5,64'h26a44f86dc13ebf8,64'hb4f484b97ef2287c,
64'haa33c7080e17a21c,64'h8fd00993ca1d8b6e,64'h6f17836eba843a91,64'hb6958c3d2b06dbd0,
64'h5e373105f57d4f1e,64'h6ed0b3601615d15b,64'h633d6bae22e5f679,64'hfffffff700080009,
64'h78d1c76d45e61927,64'h794ddd5c08f8a841,64'h07046ea6728644ae,64'he8153aa28fa6f37e,
64'h820421c9d66a62ad,64'hd70aaa2719845595,64'h19d27f3b9fd64ae7,64'h6fe9293b3c0f7e0c,
64'h1dd39fd932821f72,64'h1262ffb649f59c7f,64'h2a21e9a5a7622f92,64'h91f465c2289d10c3,
64'hedf6d2425bbc2678,64'h6a98e8187dd42b3b,64'h6ee0aa74c8022c92,64'h1fffffffe0000000,
64'hf0b4dd4c43307b04,64'h384bf401f1e761a9,64'hbf96468a8ea75ff9,64'h06f781d38d73e956,
64'h40147bf2c9fb1a97,64'hb8ca0a51b9ae9d22,64'h35227c37e09f5fbf,64'ha7a425d0f79143db,
64'h519e384570bd10db,64'h7e804ca250ec5b6c,64'h78bc1b78d421d485,64'hb4ac61ee5836de7b,
64'hf1b98831abea78ee,64'h76859b03b0ae8ad5,64'h19eb5d74172fb3c5,64'hffffffbf00400041,
64'hc68e3b6d2f30c935,64'hca6eeae347c54205,64'h3823753394322570,64'h40a9d51b7d379be9,
64'h10210e52b3531564,64'hb855513ecc22aca2,64'hce93f9dcfeb25738,64'h7f4949dce07bf05d,
64'hee9cfec99410fb90,64'h9317fdb24face3f8,64'h510f4d2e3b117c8f,64'h8fa32e1544e88614,
64'h6fb69219dde133b9,64'h54c740c6eea159d5,64'h770553a94011648d,64'hffffffff00000000,
64'h85a6ea691983d819,64'hc25fa0108f3b0d47,64'hfcb23459753affc3,64'h37bc0e9c6b9f4ab0,
64'h00a3df984fd8d4b6,64'hc6505292cd74e90b,64'ha913e1c004fafdf7,64'h3d212e8cbc8a1ed3,
64'h8cf1c22d85e886d6,64'hf40265158762db5d,64'hc5e0dbc9a10ea425,64'ha5630f77c1b6f3d3,
64'h8dcc41945f53c769,64'hb42cd820857456a5,64'hcf5aeba0b97d9e28,64'hfffffdff02000201,
64'h3471db6f798649a2,64'h537757203e2a1022,64'hc11ba99da1912b7f,64'h054ea8dde9bcdf46,
64'h810872959a98ab20,64'hc2aa89fb6115650b,64'h749fceedf592b9ba,64'hfa4a4eea03df82e5,
64'h74e7f653a087dc79,64'h98bfed967d671fbc,64'h887a6973d88be476,64'h7d1970ae2744309c,
64'h7db490d1ef099dc5,64'ha63a0639750acea6,64'hb82a9d4d008b2465,64'hfffffffefffffff9,
64'h2d37534ccc1ec0c4,64'h12fd008a79d86a32,64'he591a2d2a9d7fe11,64'hbde074e45cfa557f,
64'h051efcc27ec6a5b0,64'h3282949c6ba74852,64'h489f0e0527d7efb3,64'he9097466e450f697,
64'h678e11702f4436ac,64'ha01328b33b16dae1,64'h2f06de5308752122,64'h2b187bc30db79e93,
64'h6e620ca6fa9e3b44,64'ha166c1092ba2b523,64'h7ad75d0bcbecf13a,64'hffffefff10001001,
64'ha38edb7ccc324d0f,64'h9bbab903f150810e,64'h08dd4cf30c895bf2,64'h2a7546ef4de6fa30,
64'h084394b0d4c558fc,64'h15544fe108ab2852,64'ha4fe7772ac95cdcd,64'hd25277571efc1721,
64'ha73fb2a0043ee3c5,64'hc5ff6cb7eb38fddc,64'h43d34ba2c45f23ac,64'he8cb85743a2184dd,
64'heda48692784cee25,64'h31d031d0a856752b,64'hc154ea6d04592323,64'hfffffffeffffffc1,
64'h69ba9a6760f6061f,64'h97e80453cec35190,64'h2c8d169c4ebff081,64'hef03a727e7d2abf3,
64'h28f7e613f6352d80,64'h9414a4e45d3a428f,64'h44f8702b3ebf7d96,64'h484ba33e2287b4b1,
64'h3c708b847a21b55d,64'h0099459ed8b6d703,64'h7836f29943a9090f,64'h58c3de196dbcf497,
64'h7310653ad4f1da1d,64'h0b36084e5d15a913,64'hd6bae8615f6789cd,64'hffff7fff80008001,
64'h1c76dbeb61926873,64'hddd5c8238a84086c,64'h46ea6798644adf90,64'h53aa377b6f37d17f,
64'h421ca586a62ac7e0,64'haaa27f0845594290,64'h27f3bb9a64ae6e63,64'h9293babef7e0b902,
64'h39fd950521f71e23,64'h2ffb65c559c7eeda,64'h1e9a5d1822f91d5e,64'h465c2ba8d10c26e1,
64'h6d24349ac2677121,64'h8e818e8642b3a957,64'h0aa7536e22c91912,64'hfffffffefffffe01,
64'h4dd4d33e07b030f5,64'hbf4022a2761a8c7c,64'h6468b4e375ff8407,64'h781d39463e955f91,
64'h47bf30a0b1a96bff,64'ha0a52726e9d21474,64'h27c3815bf5fbecae,64'h425d19f3143da586,
64'he3845c24d10daae7,64'h04ca2cf6c5b6b818,64'hc1b794cd1d484875,64'hc61ef0cd6de7a4b6,
64'h988329d9a78ed0e5,64'h59b04272e8ad4898,64'hb5d74310fb3c4e62,64'hfffc000300040001,
64'he3b6df5b0c934398,64'heeae41225420435a,64'h37533cc52256fc7e,64'h9d51bbdd79be8bf6,
64'h10e52c3731563efe,64'h5513f8472aca147b,64'h3f9ddcd425737317,64'h949dd5fbbf05c80c,
64'hcfeca82a0fb8f117,64'h7fdb2e2bce3f76cf,64'hf4d2e8c117c8eaf0,64'h32e15d4888613706,
64'h6921a4d9133b8905,64'h740c7436159d4ab4,64'h553a9b711648c890,64'hfffffffefffff001,
64'h6ea699f23d8187a6,64'hfa011518b0d463db,64'h2345a71eaffc2035,64'hc0e9ca34f4aafc85,
64'h3df985078d4b5ff6,64'h0529393c4e90a39b,64'h3e1c0ae0afdf656f,64'h12e8cf9aa1ed2c2e,
64'h1c22e12d886d5731,64'h265167b62db5c0c0,64'h0dbca66eea4243a2,64'h30f786716f3d25aa,
64'hc4194ed13c768724,64'hcd821399456a44be,64'haeba188cd9e2730b,64'hffe0001f00200001,
64'h1db6fadf649a1cb9,64'h75720919a1021ac9,64'hba99e62a12b7e3ef,64'hea8ddeefcdf45fac,
64'h872961b98ab1f7f0,64'ha89fc23b5650a3d6,64'hfceee6a22b9b98b7,64'ha4eeafe1f82e405c,
64'h7f6541567dc788b2,64'hfed9716171fbb675,64'ha697460fbe475779,64'h970aea454309b82f,
64'h490d26cb99dc4825,64'ha063a1b3acea559d,64'ha9d4db8ab246447e,64'hfffffffeffff8001,
64'h7534cf94ec0c3d2d,64'hd008a8cc86a31ed1,64'h1a2d38f67fe101a7,64'h074e51ada557e422,
64'hefcc283d6a5affaf,64'h2949c9e274851cd8,64'hf0e057067efb2b77,64'h97467cd50f696170,
64'he117096c436ab988,64'h328b3db26dae05ff,64'h6de5337752121d10,64'h87bc338c79e92d4f,
64'h20ca768fe3b4391a,64'h6c109cd02b5225ea,64'h75d0c46bcf139853,64'hff0000ff01000001,
64'hedb7d6fb24d0e5c8,64'hab9048d00810d645,64'hd4cf315595bf1f73,64'h546ef7856fa2fd59,
64'h394b0dd0558fbf7c,64'h44fe11dfb2851eab,64'he77735185cdcc5b1,64'h27757f14c17202db,
64'hfb2a0ab6ee3c458d,64'hf6cb8b128fddb3a1,64'h34ba3082f23abbc3,64'hb857522e184dc174,
64'h4869365ecee24126,64'h031d0da26752ace3,64'h4ea6dc5a923223eb,64'hfffffffefffc0001,
64'ha9a67caa6061e965,64'h8045466a3518f682,64'hd169c7b3ff080d38,64'h3a728d6d2abf2110,
64'h7e6141f252d7fd71,64'h4a4e4f14a428e6bf,64'h8702b83af7d95bb1,64'hba33e6ac7b4b0b7c,
64'h08b84b691b55cc39,64'h9459ed946d702ff7,64'h6f299bbd9090e87d,64'h3de19c67cf496a74,
64'h0653b4801da1c8cf,64'h6084e6845a912f4d,64'hae862361789cc295,64'hf80007ff08000001,
64'h6dbeb7e026872e39,64'h5c8246854086b223,64'ha6798ab2adf8fb92,64'ha377bc2d7d17eac6,
64'hca586e83ac7dfbdf,64'h27f08eff9428f556,64'h3bb9a8c9e6e62d81,64'h3babf8a70b9016d7,
64'hd95055be71e22c61,64'hb65c589b7eed9d01,64'ha5d1841891d5de17,64'hc2ba9175c26e0b9b,
64'h4349b2f87712092e,64'h18e86d133a956718,64'h7536e2d691911f56,64'hfffffffeffe00001,
64'h4d33e558030f4b23,64'h022a3355a8c7b40c,64'h8b4e3da5f84069ba,64'hd3946b6a55f9087f,
64'hf30a0f9596bfeb85,64'h527278a7214735f6,64'h3815c1dbbecadd84,64'hd19f3568da585bdb,
64'h45c25b48daae61c8,64'ha2cf6ca76b817fb4,64'h794cddef848743e5,64'hef0ce33f7a4b539f,
64'h329da400ed0e4678,64'h04273425d4897a65,64'h74311b10c4e614a3,64'hc0003fff40000001,
64'h6df5bf04343971c5,64'he412342c04359116,64'h33cc559a6fc7dc8b,64'h1bbde170e8bf562b,
64'h52c3742363efdef2,64'h3f8477fda147aaaf,64'hddcd465037316c07,64'hdd5fc5395c80b6b7,
64'hca82adf98f116302,64'hb2e2c4e0f76ce803,64'h2e8c20c98eaef0b3,64'h15d48bb413705cd2,
64'h1a4d97c5b890496e,64'hc7436899d4ab38c0,64'ha9b716b78c88faad,64'hfffffffeff000001,
64'h699f2ac2187a5916,64'h11519aad463da060,64'h5a71ed33c2034dcc,64'h9ca35b58afc843f2,
64'h98507cb3b5ff5c21,64'h9393c53b0a39afae,64'hc0ae0edef656ec1f,64'h8cf9ab4cd2c2ded2,
64'h2e12da48d5730e3e,64'h167b65405c0bfd9b,64'hca66ef7f243a1f25,64'h78671a02d25a9cf1,
64'h94ed2008687233bf,64'h2139a12ea44bd328,64'ha188d8892730a515,64'h0002000000000002,
64'h6fadf824a1cb8e25,64'h2091a16721ac88a9,64'h9e62acd47e3ee457,64'hddef0b8745fab158,
64'h961ba11d1f7ef78e,64'hfc23bfee0a3d5577,64'hee6a3287b98b6032,64'heafe29d0e405b5b2,
64'h54156fd2788b180a,64'h9716270cbb674013,64'h7461064d75778597,64'haea45da09b82e690,
64'hd26cbe2dc4824b70,64'h3a1b44d4a559c5fa,64'h4db8b5c16447d563,64'hfffffffef8000001,
64'h4cf95613c3d2c8ad,64'h8a8cd56a31ed0300,64'hd38f69a0101a6e5e,64'he51adac97e421f8c,
64'hc283e5a1affae104,64'h9c9e29dc51cd7d6c,64'h057076fdb2b760f2,64'h67cd5a6a9616f68c,
64'h7096d247ab9871ef,64'hb3db2a02e05fecd8,64'h53377bff21d0f922,64'hc338d01992d4e785,
64'ha769004743919df4,64'h09cd0976225e993f,64'h0c46c44e398528a3,64'h0010000000000010,
64'h7d6fc1280e5c7125,64'h048d0b3a0d644547,64'hf31566a7f1f722b4,64'hef785c402fd58aba,
64'hb0dd08ecfbf7bc6c,64'he11dff7751eaabb1,64'h73519444cc5b0189,64'h57f14e8e202dad89,
64'ha0ab7e95c458c04e,64'hb8b13869db3a0094,64'ha308326eabbc2cb5,64'h7522ed09dc17347b,
64'h9365f17424125b7a,64'hd0da26a62ace2fcf,64'h6dc5ae0d223eab16,64'hfffffffec0000001,
64'h67cab0a01e964566,64'h5466ab558f6817fc,64'h9c7b4d0680d372ea,64'h28d6d652f210fc59,
64'h141f2d137fd7081a,64'he4f14ee68e6beb5c,64'h2b83b7ed95bb0790,64'h3e6ad357b0b7b45d,
64'h84b692405cc38f75,64'h9ed9501c02ff66bb,64'h99bbdffb0e87c90e,64'h19c680d296a73c22,
64'h3b48023f1c8cef9b,64'h4e684bb112f4c9f8,64'h62362271cc294518,64'h0080000000000080,
64'heb7e094372e38925,64'h246859d06b222a38,64'h98ab35468fb91599,64'h7bc2e2087eac55c9,
64'h86e8476cdfbde35b,64'h08effbc18f555d81,64'h9a8ca22962d80c45,64'hbf8a7473016d6c46,
64'h055bf4b322c6026b,64'hc589c353d9d0049b,64'h1841937a5de165a3,64'ha9176851e0b9a3d5,
64'h9b2f8ba52092dbcc,64'h86d1353756717e72,64'h6e2d706c11f558ad,64'hfffffffd00000001,
64'h3e558503f4b22b2d,64'ha3355aae7b40bfde,64'he3da6838069b974c,64'h46b6b2989087e2c7,
64'ha0f9689bfeb840d0,64'h278a773b735f5ad9,64'h5c1dbf6dadd83c7f,64'hf3569abe85bda2e7,
64'h25b49206e61c7ba4,64'hf6ca80e417fb35d4,64'hcddeffdc743e486c,64'hce340694b539e110,
64'hda4011f9e4677cd7,64'h73425d8a97a64fbe,64'h11b11391614a28bd,64'h0400000000000400,
64'h5bf04a22971c4921,64'h2342ce84591151bf,64'hc559aa387dc8acc4,64'hde171046f562ae45,
64'h37423b6afdef1ad4,64'h477fde0c7aaaec08,64'hd465114f16c06224,64'hfc53a39d0b6b622b,
64'h2adfa59916301358,64'h2c4e1aa4ce8024d2,64'hc20c9bd2ef0b2d18,64'h48bb429405cd1ea3,
64'hd97c5d2d0496de5c,64'h3689a9beb38bf38c,64'h716b83638faac565,64'hffffffef00000001,
64'hf2ac2820a5915967,64'h19aad578da05feeb,64'h1ed341c734dcba59,64'h35b594c6843f1636,
64'h07cb44e4f5c2067b,64'h3c53b9dc9afad6c7,64'he0edfb6f6ec1e3f6,64'h9ab4d5fb2ded1731,
64'h2da4903830e3dd1f,64'hb6540727bfd9ae99,64'h6ef7fee9a1f2435a,64'h71a034aba9cf087a,
64'hd2008fd5233be6b2,64'h9a12ec57bd327ded,64'h8d889c8b0a5145e8,64'h2000000000002000,
64'hdf825116b8e24906,64'h1a167423c88a8df7,64'h2acd51c9ee45661a,64'hf0b8823dab157222,
64'hba11db58ef78d69f,64'h3bfef065d557603e,64'ha3288a7eb603111a,64'he29d1cef5b5b1151,
64'h56fd2cc9b1809abf,64'h6270d5277401268f,64'h1064de9d785968ba,64'h45da14a22e68f516,
64'hcbe2e96e24b6f2da,64'hb44d4df69c5f9c5f,64'h8b5c1b1f7d562b25,64'hffffff7f00000001,
64'h9561410c2c8acb31,64'hcd56abc6d02ff758,64'hf69a0e39a6e5d2c8,64'hadaca63521f8b1af,
64'h3e5a2727ae1033d8,64'he29dcee5d7d6b637,64'h076fdb82760f1fa9,64'hd5a6afdd6f68b984,
64'h6d2481c2871ee8f7,64'hb2a03942fecd74c3,64'h77bff7500f921acd,64'h8d01a5604e7843cd,
64'h90047eaf19df358a,64'hd09762c1e993ef64,64'h6c44e45c528a2f3c,64'h000000010000ffff,
64'hfc1288bbc712482a,64'hd0b3a11e44546fb8,64'h566a8e50722b30cf,64'h85c411f458ab9109,
64'hd08edacc7bc6b4f3,64'hdff7832faabb01ef,64'h194453fab01888cb,64'h14e8e781dad88a81,
64'hb7e9664f8c04d5f6,64'h1386a93ea0093475,64'h8326f4ebc2cb45d0,64'h2ed0a5137347a8ae,
64'h5f174b7725b796ca,64'ha26a6fb9e2fce2f3,64'h5ae0d8ffeab15924,64'hfffffbff00000001,
64'hab0a086564565984,64'h6ab55e3c817fbaba,64'hb4d071d4372e9639,64'h6d6531ae0fc58d73,
64'hf2d1393e70819ebf,64'h14ee7735beb5b1b1,64'h3b7edc13b078fd48,64'had357ef17b45cc1a,
64'h69240e1738f747b5,64'h9501ca1cf66ba613,64'hbdffba837c90d665,64'h680d2b0673c21e64,
64'h8023f57ccef9ac4c,64'h84bb16154c9f7b1a,64'h622722e5945179dd,64'h000000080007fff8,
64'he09445e538924149,64'h859d08f822a37dba,64'hb354728591598676,64'h2e208fa6c55c8844,
64'h8476d669de35a792,64'hffbc198355d80f72,64'hca229fd580c44658,64'ha7473c0ed6c45408,
64'hbf4b32816026afab,64'h9c3549f50049a3a8,64'h1937a762165a2e7c,64'h7685289c9a3d456f,
64'hf8ba5bbb2dbcb64e,64'h13537dd417e71793,64'hd706c801558ac91e,64'hffffdfff00000001,
64'h5850433022b2cc1b,64'h55aaf1e70bfdd5cd,64'ha6838ea6b974b1c3,64'h6b298d737e2c6b95,
64'h9689c9fa840cf5f1,64'ha773b9adf5ad8d88,64'hdbf6e09e83c7ea3f,64'h69abf790da2e60cb,
64'h492070bcc7ba3da5,64'ha80e50ebb35d3094,64'heffdd420e486b323,64'h406958369e10f31d,
64'h011fabea77cd625c,64'h25d8b0ae64fbd8cc,64'h1139172fa28bcee5,64'h00000040003fffc0,
64'h04a22f30c4920a41,64'h2ce847c5151bedcc,64'h9aa394318acc33ab,64'h71047d372ae4421f,
64'h23b6b352f1ad3c8c,64'hfde0cc21aec07b89,64'h5114feb2062232ba,64'h3a39e07bb622a03b,
64'hfa59941001357d53,64'he1aa4fac024d1d3c,64'hc9bd3b10b2d173e0,64'hb42944e7d1ea2b75,
64'hc5d2dde06de5b269,64'h9a9beea0bf38bc98,64'hb8364010ac5648ea,64'hfffeffff00000001,
64'hc2821983159660d6,64'had578f3a5feeae66,64'h341c753acba58e13,64'h594c6b9ef1635ca5,
64'hb44e4fd82067af84,64'h3b9dcd74ad6c6c3b,64'hdfb704fa1e3f51f2,64'h4d5fbc89d1730655,
64'h490385e83dd1ed26,64'h407287629ae9849b,64'h7feea10e24359911,64'h034ac1b6f08798e6,
64'h08fd5f53be6b12e0,64'h2ec5857427dec65f,64'h89c8b97d145e7728,64'h0000020001fffe00,
64'h2511798624905208,64'h67423e29a8df6e5f,64'hd51ca19056619d54,64'h8823e9bc572210f5,
64'h1db59a988d69e45f,64'hef0661147603dc41,64'h88a7f592311195ce,64'hd1cf03deb11501d7,
64'hd2cca08709abea91,64'h0d527d671268e9d9,64'h4de9d88b968b9efa,64'ha14a27438f515ba3,
64'h2e96ef096f2d9342,64'hd4df7509f9c5e4bc,64'hc1b2008a62b2474b,64'hfff7ffff00000001,
64'h1410cc1eacb306aa,64'h6abc79d7ff75732b,64'ha0e3a9d75d2c7097,64'hca635cf98b1ae526,
64'ha2727ec6033d7c1b,64'hdcee6ba66b6361d7,64'hfdb827d6f1fa8f8a,64'h6afde4508b9832a6,
64'h481c2f43ee8f692e,64'h03943b16d74c24d6,64'hff75087421acc885,64'h1a560db7843cc730,
64'h47eafa9df3589700,64'h762c2ba23ef632f7,64'h4e45cbeca2f3b93c,64'h000010000ffff000,
64'h288bcc322482903f,64'h3a11f15046fb72f5,64'ha8e50c88b30cea9a,64'h411f4de6b91087a4,
64'hedacd4c46b4f22f8,64'h783308aab01ee201,64'h453fac95888cae6c,64'h8e781efb88a80eb2,
64'h9665043e4d5f5482,64'h6a93eb3893474ec8,64'h6f4ec45eb45cf7ce,64'h0a513a217a8add13,
64'h74b7784c796c9a0f,64'ha6fba855ce2f25da,64'h0d90045915923a52,64'hffbfffff00000001,
64'ha08660f565983550,64'h55e3cec2fbab9955,64'h071d4ebfe96384b3,64'h531ae7d258d7292a,
64'h1393f63519ebe0d3,64'he7735d395b1b0eb2,64'hedc13ebe8fd47c49,64'h57ef22875cc1952d,
64'h40e17a21747b496e,64'h1ca1d8b6ba6126b0,64'hfba843a80d664421,64'hd2b06dbc21e63980,
64'h3f57d4f19ac4b7fe,64'hb1615d14f7b197b5,64'h722e5f67179dc9de,64'h000080007fff8000,
64'h445e6192241481f7,64'hd08f8a8337db97a7,64'h4728644a986754cb,64'h08fa6f37c8843d1e,
64'h6d66a62a5a7917b9,64'hc198455880f71005,64'h29fd64ae4465735e,64'h73c0f7e04540758c,
64'hb32821f66afaa40c,64'h549f59c79a3a763d,64'h7a7622f8a2e7be6d,64'h5289d10bd456e898,
64'ha5bbc266cb64d075,64'h37dd42b371792ecb,64'h6c8022c8ac91d290,64'hfdffffff00000001,
64'h043307b02cc1aa7b,64'haf1e7619dd5ccaa6,64'h38ea75ff4b1c2598,64'h98d73e94c6b9494e,
64'h9c9fb1a8cf5f0698,64'h3b9ae9d1d8d87589,64'h6e09f5fb7ea3e241,64'hbf79143ce60ca966,
64'h070bd10da3da4b6e,64'he50ec5b5d3093580,64'hdd421d476b322101,64'h95836de70f31cbfa,
64'hfabea78dd625bfef,64'h8b0ae8acbd8cbda3,64'h9172fb3bbcee4eed,64'h00040003fffc0000,
64'h22f30c9320a40fb6,64'h847c541fbedcbd32,64'h39432256c33aa656,64'h47d379be4421e8f0,
64'h6b353155d3c8bdc5,64'h0cc22aca07b88022,64'h4feb2573232b9aef,64'h9e07bf052a03ac5d,
64'h99410fb857d5205b,64'ha4face3ed1d3b1e6,64'hd3b117c8173df365,64'h944e8860a2b744be,
64'h2dde133b5b2683a3,64'hbeea159c8bc97657,64'h64011648648e947d,64'hefffffff00000001,
64'h21983d81660d53d8,64'h78f3b0d3eae6552b,64'hc753affb58e12cbf,64'hc6b9f4aa35ca4a6c,
64'he4fd8d4a7af834bc,64'hdcd74e8fc6c3ac47,64'h704fafdef51f1205,64'hfbc8a1ec30654b2b,
64'h385e886d1ed25b70,64'h28762db59849abf9,64'hea10ea4159910802,64'hac1b6f3c798e5fcc,
64'hd5f53c75b12dff71,64'h58574569ec65ed14,64'h8b97d9e1e7727764,64'h0020001fffe00000,
64'h1798649a05207daf,64'h23e2a101f6e5e98c,64'hca1912b719d532af,64'h3e9bcdf4210f477e,
64'h59a98ab19e45ee25,64'h661156503dc40110,64'h7f592b9b195cd776,64'hf03df82d501d62e4,
64'hca087dc6bea902d4,64'h27d671fb8e9d8f2b,64'h9d88be46b9ef9b22,64'ha274430915ba25ec,
64'h6ef099dbd9341d17,64'hf750ace95e4bb2b3,64'h2008b2462474a3e5,64'h7fffffff00000001,
64'h0cc1ec0c306a9ebf,64'hc79d86a25732a955,64'h3a9d7fe0c70965f2,64'h35cfa557ae52535a,
64'h27ec6a5ad7c1a5d9,64'he6ba7484361d6232,64'h827d7efaa8f89025,64'hde450f68832a5951,
64'hc2f44369f692db7f,64'h43b16dadc24d5fc7,64'h50875211cc884009,64'h60db79e8cc72fe5b,
64'hafa9e3b3896ffb82,64'hc2ba2b51632f689e,64'h5cbecf133b93bb1c,64'h010000ffff000000,
64'hbcc324d02903ed78,64'h1f150810b72f4c5f,64'h50c895becea99572,64'hf4de6fa2087a3bef,
64'hcd4c558ef22f7126,64'h308ab284ee20087d,64'hfac95cdbcae6bbad,64'h81efc17180eb1719,
64'h5043ee3bf548169a,64'h3eb38fdd74ec7957,64'hec45f239cf7cd90c,64'h13a2184dadd12f5b,
64'h7784cee1c9a0e8b5,64'hba856751f25d9591,64'h0045923223a51f27,64'hfffffffb00000005,
64'h660f60618354f5f8,64'h3cec3518b9954aa2,64'hd4ebff07384b2f8f,64'hae7d2abe72929acf,
64'h3f6352d7be0d2ec7,64'h35d3a428b0eb1189,64'h13ebf7d947c48124,64'hf2287b4a1952ca82,
64'h17a21b55b496dbf2,64'h1d8b6d70126afe36,64'h843a909064420046,64'h06dbcf496397f2d5,
64'h7d4f1da14b7fdc0b,64'h15d15a91197b44ea,64'he5f6789bdc9dd8de,64'h080007fff8000000,
64'he6192686481f6bbb,64'hf8a84085b97a62f8,64'h8644adf8754cab8e,64'ha6f37d1743d1df71,
64'h6a62ac7d917b892a,64'h84559428710043e7,64'hd64ae6e55735dd61,64'h0f7e0b900758b8c4,
64'h821f71e1aa40b4ce,64'hf59c7eeca763cab7,64'h622f91d57be6c859,64'h9d10c26d6e897ad8,
64'hbc2677114d0745a5,64'hd42b3a9492ecac83,64'h022c91911d28f938,64'hffffffdf00000021,
64'h307b030f1aa7afbd,64'he761a8c6ccaa550f,64'ha75ff83fc2597c72,64'h73e955f89494d673,
64'hfb1a96bef0697637,64'hae9d214687588c47,64'h9f5fbeca3e240920,64'h9143da57ca965409,
64'hbd10daada4b6df90,64'hec5b6b809357f1b0,64'h21d484872210022c,64'h36de7a4b1cbf96a8,
64'hea78ed0d5bfee055,64'hae8ad488cbda2750,64'h2fb3c4e5e4eec6e9,64'h40003fffc0000000,
64'h30c9343940fb5dd1,64'hc5420434cbd317b9,64'h32256fc7aa655c6c,64'h379be8bf1e8efb83,
64'h531563ef8bdc494d,64'h22aca14788021f34,64'hb2573730b9aeeb02,64'h7bf05c803ac5c620,
64'h10fb8f115205a66c,64'hace3f76c3b1e55b1,64'h117c8eaedf3642c5,64'he886136f744bd6bc,
64'he133b88f683a2d23,64'ha159d4aa97656412,64'h11648c88e947c9c0,64'hfffffeff00000101,
64'h83d81879d53d7de7,64'h3b0d463d6552a871,64'h3affc20312cbe38b,64'h9f4aafc7a4a6b395,
64'hd8d4b5fe834bb1b1,64'h74e90a393ac46233,64'hfafdf655f12048fc,64'h8a1ed2c254b2a044,
64'he886d57225b6fc7b,64'h62db5c0b9abf8d79,64'h0ea4243a1080115f,64'hb6f3d259e5fcb53f,
64'h53c76871dff702a1,64'h7456a44b5ed13a7b,64'h7d9e273027763747,64'h0001fffffffffffe,
64'h8649a1cb07daee87,64'h2a1021ac5e98bdc2,64'h912b7e3e532ae35f,64'hbcdf45f9f477dc17,
64'h98ab1f7e5ee24a66,64'h15650a3d4010f99f,64'h92b9b98acd77580b,64'hdf82e404d62e30fd,
64'h87dc788a902d3360,64'h671fbb66d8f2ad83,64'h8be47576f9b21628,64'h44309b82a25eb5d9,
64'h099dc48241d16911,64'h0acea559bb2b208b,64'h8b2464474a3e4e00,64'hfffff7ff00000801,
64'h1ec0c3d2a9ebef34,64'hd86a31ec2a954387,64'hd7fe1019965f1c57,64'hfa557e4125359ca4,
64'hc6a5affa1a5d8d82,64'ha74851ccd6231195,64'hd7efb2b6890247d9,64'h50f69616a595021c,
64'h4436ab982db7e3d1,64'h16dae05fd5fc6bc5,64'h752121d084008af8,64'hb79e92d42fe5a9f3,
64'h9e3b4390ffb81506,64'ha2b5225df689d3d5,64'hecf139843bb1ba35,64'h000ffffffffffff0,
64'h324d0e5c3ed77434,64'h50810d63f4c5ee0f,64'h895bf1f699571af4,64'he6fa2fd4a3bee0b3,
64'hc558fbf6f712532c,64'hab2851ea0087ccf8,64'h95cdcc5a6bbac054,64'hfc17202cb17187e2,
64'h3ee3c45881699afc,64'h38fddb39c7956c15,64'h5f23abbbcd90b13c,64'h2184dc1712f5aec6,
64'h4cee24120e8b4888,64'h56752acdd9590458,64'h5923223e51f26ffc,64'hffffbfff00004001,
64'hf6061e954f5f79a0,64'hc3518f6754aa1c32,64'hbff080d2b2f8e2b2,64'hd2abf21029ace519,
64'h352d7fd6d2ec6c0a,64'h3a428e6bb1188ca3,64'hbf7d95ba48123ec2,64'h87b4b0b72ca810de,
64'h21b55cc36dbf1e86,64'hb6d702feafe35e28,64'ha9090e87200457bd,64'hbcf496a67f2d4f93,
64'hf1da1c8bfdc0a82c,64'h15a912f4b44e9ea3,64'h6789cc28dd8dd1a1,64'h007fffffffffff80,
64'h926872e2f6bba19f,64'h84086b21a62f7076,64'h4adf8fb8cab8d79c,64'h37d17eac1df70591,
64'h2ac7dfbdb892995a,64'h59428f55043e67bb,64'hae6e62d75dd6029c,64'he0b9016c8b8c3f09,
64'hf71e22c50b4cd7df,64'hc7eed9cf3cab60a7,64'hf91d5de06c8589de,64'h0c26e0b997ad762f,
64'h67712092745a443e,64'hb3a95670cac822be,64'hc91911f48f937fde,64'hfffdffff00020001,
64'hb030f4b17afbccf9,64'h1a8c7b40a550e18a,64'hff84069a97c7158b,64'h955f90874d6728c2,
64'ha96bfeb79763604f,64'hd214735e88c46517,64'hfbecadd74091f60b,64'h3da585bd654086ec,
64'h0daae61c6df8f42f,64'hb6b817fa7f1af13b,64'h4848743e0022bde3,64'he7a4b538f96a7c93,
64'h8ed0e466ee054159,64'had4897a5a274f518,64'h3c4e6149ec6e8d05,64'h03fffffffffffc00,
64'h9343971bb5dd0cf4,64'h20435911317b83ac,64'h56fc7dc855c6bcde,64'hbe8bf561efb82c87,
64'h563efdeec494cacf,64'hca147aaa21f33dd6,64'h737316bfeeb014db,64'h05c80b6b5c61f841,
64'hb8f1162f5a66bef1,64'h3f76ce7fe55b0532,64'hc8eaef0a642c4ee9,64'h613705ccbd6bb178,
64'h3b890496a2d221ed,64'h9d4ab38b564115eb,64'h48c88faa7c9bfeea,64'hffefffff00100001,
64'h8187a590d7de67c3,64'hd463da052a870c50,64'hfc2034dbbe38ac51,64'haafc843e6b39460c,
64'h4b5ff5c1bb1b0273,64'h90a39afa462328b2,64'hdf656ec1048fb051,64'hed2c2dec2a04375f,
64'h6d5730e36fc7a178,64'hb5c0bfd8f8d789d3,64'h4243a1f20115ef16,64'h3d25a9cecb53e491,
64'h7687233b702a0ac4,64'h6a44bd3213a7a8bb,64'he2730a5063746827,64'h1fffffffffffe000,
64'h9a1cb8e1aee8679c,64'h021ac88a8bdc1d5f,64'hb7e3ee44ae35e6ee,64'hf45fab147dc16433,
64'hb1f7ef7824a65676,64'h50a3d5570f99eeaa,64'h9b98b6027580a6d5,64'h2e405b5ae30fc208,
64'hc788b17fd335f783,64'hfbb674002ad8298f,64'h4757785921627742,64'h09b82e68eb5d8bbd,
64'hdc4824b616910f67,64'hea559c5eb208af54,64'h46447d55e4dff74e,64'hff7fffff00800001,
64'h0c3d2c8abef33e14,64'ha31ed02f5438627a,64'he101a6e4f1c56281,64'h57e421f859ca305b,
64'h5affae0fd8d81396,64'h851cd7d63119458c,64'hfb2b760e247d8282,64'h69616f685021baf1,
64'h6ab9871e7e3d0bbd,64'hae05feccc6bc4e93,64'h121d0f9208af78ae,64'he92d4e775a9f2487,
64'hb43919de8150561d,64'h5225e9939d3d45d5,64'h1398528a1ba34131,64'h00000000fffeffff,
64'hd0e5c71177433cdc,64'h10d644545ee0eaf8,64'hbf1f722a71af376b,64'ha2fd58aaee0b2191,
64'h8fbf7bc62532b3ab,64'h851eaaba7ccf754e,64'hdcc5b017ac0536a4,64'h7202dad8187e103f,
64'h3c458c0499afbc12,64'hddb3a00856c14c71,64'h3abbc2cb0b13ba0e,64'h4dc173475aec5de8,
64'he24125b6b4887b32,64'h52ace2fc90457a99,64'h3223eab126ffba6e,64'hfbffffff04000001,
64'h61e96455f799f0a0,64'h18f6817fa1c313cb,64'h080d372e8e2b1401,64'hbf210fc4ce5182d6,
64'hd7fd7080c6c09cae,64'h28e6beb588ca2c5c,64'hd95bb07823ec1409,64'h4b0b7b45810dd785,
64'h55cc38f6f1e85de5,64'h702ff66b35e27493,64'h90e87c90457bc570,64'h496a73c1d4f92431,
64'ha1c8cef90a82b0e3,64'h912f4c9ee9ea2ea6,64'h9cc29450dd1a0988,64'h00000007fff7fff8,
64'h872e3891ba19e6da,64'h86b222a2f70757c0,64'hf8fb91588d79bb53,64'h17eac55c70590c83,
64'h7dfbde3529959d54,64'h28f555d7e67baa6c,64'he62d80c36029b51a,64'h9016d6c3c3f081f5,
64'he22c6025cd7de08f,64'hed9d0048b60a6382,64'hd5de1659589dd06f,64'h6e0b9a3cd762ef3e,
64'h12092dbca443d989,64'h956717e6822bd4c6,64'h911f558a37fdd36f,64'hdfffffff20000001,
64'h0f4b22b2bccf84fd,64'hc7b40bfd0e189e58,64'h4069b9747158a008,64'hf9087e2b728c16ab,
64'hbfeb840c3604e56a,64'h4735f5ad465162df,64'hcadd83c71f60a042,64'h585bda2e086ebc26,
64'hae61c7b98f42ef26,64'h817fb35caf13a495,64'h8743e4862bde2b7c,64'h4b539e10a7c92186,
64'h0e4677cd54158713,64'h897a64fb4f51752c,64'he614a28ae8d04c3c,64'h0000003fffbfffc0,
64'h3971c491d0cf36cc,64'h3591151bb83abdfc,64'hc7dc8acb6bcdda91,64'hbf562ae382c86418,
64'hefdef1ac4cacea9d,64'h47aaaec033dd535f,64'h316c0622014da8c9,64'h80b6b6221f840fa4,
64'h116301356bef0471,64'h6ce8024cb0531c09,64'haef0b2d0c4ee8372,64'h705cd1e9bb1779ed,
64'h90496de5221ecc48,64'hab38bf38115ea62c,64'h88faac55bfee9b74,64'h0000000000000001
};
  //------------------------
  // 512
  //------------------------
  localparam [2*512-1:0][63:0] NTT_GF64_BWD_N512_PHI_L = {
64'h3da05fee70c4f2ba,64'hc843f1629460b551,64'h39afad6c328b16f6,64'hc2ded1724375e12e,
64'h0bfd9ae9789d24a4,64'h5a9cf0873e490c2e,64'h4bd327de7a8ba95c,64'h000001fffdfffe00,
64'hac88a8dec1d5efdf,64'hfab15721164320bb,64'h3d5576039eea9af6,64'h05b5b114fc207d1c,
64'h674012688298e045,64'h82e68f50d8bbcf65,64'h59c5f9c58af5315b,64'h0000000000000008,
64'hed02ff74862795cf,64'h421f8b1aa305aa82,64'hcd7d6b629458b7af,64'h16f68b981baf096a,
64'h5fecd74bc4e92520,64'hd4e7843bf248616e,64'h5e993ef5d45d4ade,64'h00000fffeffff000,
64'h644546fb0eaf7ef3,64'hd58ab90fb21905d1,64'heaabb01df754d7af,64'h2dad88a7e103e8e0,
64'h3a00934714c70225,64'h17347a8ac5de7b24,64'hce2fce2e57a98ad6,64'h0000000000000040,
64'h6817fbab313cae71,64'h10fc58d7182d540e,64'h6beb5b1aa2c5bd72,64'hb7b45cc0dd784b50,
64'hff66ba60274928fe,64'ha73c21e592430b6a,64'hf4c9f7b0a2ea56ee,64'h00007fff7fff8000,
64'h222a37db757bf795,64'hac55c88390c82e82,64'h555d80f6baa6bd71,64'h6d6c4540081f46ff,
64'hd0049a39a6381127,64'hb9a3d4562ef3d920,64'h717e7178bd4c56aa,64'h0000000000000200,
64'h40bfdd5c89e57385,64'h87e2c6b8c16aa070,64'h5f5ad8d8162deb8d,64'hbda2e60bebc25a7b,
64'hfb35d3083a4947e9,64'h39e10f3192185b4b,64'ha64fbd8c1752b769,64'h0003fffbfffc0000,
64'h1151bedcabdfbca7,64'h62ae44218641740b,64'haaec07b7d535eb86,64'h6b622a0340fa37f5,
64'h8024d1d331c08932,64'hcd1ea2b6779ec8fb,64'h8bf38bc8ea62b54d,64'h0000000000001000,
64'h05feeae64f2b9c26,64'h3f1635ca0b55037c,64'hfad6c6c2b16f5c66,64'hed1730645e12d3d3,
64'hd9ae9848d24a3f41,64'hcf08798d90c2da57,64'h327dec65ba95bb43,64'h001fffdfffe00000,
64'h8a8df6e55efde538,64'h1572210f320ba055,64'h57603dc3a9af5c2b,64'h5b11501d07d1bfa5,
64'h01268e9d8e04498c,64'h68f515b9bcf647d2,64'h5f9c5e4b5315aa64,64'h0000000000008000,
64'h2ff75732795ce130,64'hf8b1ae515aa81bdf,64'hd6b6361c8b7ae329,64'h68b98329f0969e91,
64'hcd74c24c9251fa02,64'h7843cc728616d2b2,64'h93ef632ed4adda17,64'h00fffeffff000000,
64'h546fb72ef7ef29bc,64'hab910879905d02a8,64'hbb01ee1f4d7ae156,64'hd88a80ea3e8dfd26,
64'h093474ec70224c60,64'h47a8add0e7b23e8d,64'hfce2f25c98ad531e,64'h0000000000040000,
64'h7fbab994cae7097f,64'hc58d7291d540def1,64'hb5b1b0ea5bd71942,64'h45cc195284b4f485,
64'h6ba6126a928fd00a,64'hc21e639730b6958d,64'h9f7b197aa56ed0b4,64'h07fff7fff8000000,
64'ha37db979bf794dde,64'h5c8843d182e8153b,64'hd80f70ff6bd70aab,64'hc4540757f46fe92a,
64'h49a3a76381126300,64'h3d456e893d91f466,64'he71792ebc56a98e9,64'h0000000000200000,
64'hfdd5cca957384bf5,64'h2c6b9494aa06f782,64'had8d8757deb8ca0b,64'h2e60ca9625a7a426,
64'h5d309357947e804d,64'h10f31cbf85b4ac62,64'hfbd8cbd92b76859c,64'h3fffbfffc0000000,
64'h1bedcbd2fbca6eeb,64'he4421e8e1740a9d6,64'hc07b88015eb85552,64'h22a03ac5a37f494a,
64'h4d1d3b1e089317fe,64'hea2b744aec8fa32f,64'h38bc97652b54c741,64'h0000000001000000,
64'heeae6551b9c25fa1,64'h635ca4a65037bc0f,64'h6c6c3ac3f5c65053,64'h730654b22d3d212f,
64'he9849abea3f40266,64'h8798e5fc2da56310,64'hdec65ed05bb42cd9,64'hfffdfffeffffffff,
64'hdf6e5e97de537758,64'h2210f477ba054ea9,64'h03dc4010f5c2aa8a,64'h1501d62e1bfa4a4f,
64'h68e9d8f24498bfee,64'h515ba25e647d1971,64'hc5e4bb2a5aa63a07,64'h0000000008000000,
64'h75732a94ce12fd01,64'h1ae5253581bde075,64'h6361d622ae328295,64'h9832a59469e90975,
64'h4c24d5fc1fa01329,64'h3cc72fe56d2b187c,64'hf632f688dda166c2,64'hffeffffefffffff1,
64'hfb72f4c4f29bbaba,64'h1087a3bed02a7547,64'h1ee20087ae155450,64'ha80eb170dfd25278,
64'h474ec79524c5ff6d,64'h8add12f523e8cb86,64'h2f25d958d531d032,64'h0000000040000000,
64'hab9954a97097e805,64'hd72929ac0def03a8,64'h1b0eb118719414a5,64'hc1952ca74f484ba4,
64'h6126afe2fd009946,64'he6397f2c6958c3df,64'hb197b44ded0b3609,64'hff7ffffeffffff81,
64'hdb97a62e94ddd5c9,64'h843d1df68153aa38,64'hf710043d70aaa280,64'h40758b8bfe9293bb,
64'h3a763cab262ffb66,64'h56e897ad1f465c2c,64'h792ecac7a98e818f,64'h0000000200000000,
64'h5ccaa55084bf4023,64'hb9494d666f781d3a,64'hd87588c38ca0a528,64'h0ca965407a425d1a,
64'h09357f1ae804ca2d,64'h31cbf96a4ac61ef1,64'h8cbda2746859b043,64'hfbfffffefffffc01,
64'hdcbd317aa6eeae42,64'h21e8efb80a9d51bc,64'hb88021f2855513f9,64'h03ac5c61f4949dd6,
64'hd3b1e55a317fdb2f,64'hb744bd6afa32e15e,64'hc97656404c740c75,64'h0000001000000000,
64'he6552a8625fa0116,64'hca4a6b387bc0e9cb,64'hc3ac46226505293a,64'h654b2a03d212e8d0,
64'h49abf8d740265168,64'h8e5fcb535630f787,64'h65ed13a742cd8214,64'hdffffffeffffe001,
64'he5e98bdb3775720a,64'h0f477dc154ea8ddf,64'hc4010f992aa89fc3,64'h1d62e30fa4a4eeb0,
64'h9d8f2ad78bfed972,64'hba25eb5cd1970aeb,64'h4bb2b20863a063a2,64'h0000008000000000,
64'h32a954382fd008a9,64'h525359c9de074e52,64'h1d623119282949ca,64'h2a5950219097467d,
64'h4d5fc6bc01328b3e,64'h72fe5a9eb187bc34,64'h2f689d3d166c109d,64'hfffffffdffff0002,
64'h2f4c5ee0bbab9049,64'h7a3bee0aa7546ef8,64'h20087ccf5544fe12,64'heb17187d25277580,
64'hec7956c05ff6cb8c,64'hd12f5aeb8cb85753,64'h5d9590451d031d0e,64'h0000040000000000,
64'h954aa1c27e804547,64'h929ace50f03a728e,64'heb1188c9414a4e50,64'h52ca810d84ba33e7,
64'h6afe35e2099459ee,64'h97f2d4f88c3de19d,64'h7b44e9e9b36084e7,64'hfffffff6fff80009,
64'h7a62f706dd5c8247,64'hd1df70583aa377bd,64'h0043e67baa27f08f,64'h58b8c3f0293babf9,
64'h63cab609ffb65c59,64'h897ad76265c2ba92,64'hecac822ae818e86e,64'h0000200000000000,
64'haa550e17f4022a34,64'h94d6728b81d3946c,64'h588c46510a527279,64'h9654086e25d19f36,
64'h57f1af134ca2cf6d,64'hbf96a7c861ef0ce4,64'hda274f509b042735,64'hffffffbeffc00041,
64'hd317b839eae41235,64'h8efb82c7d51bbde2,64'h021f33dd513f8478,64'hc5c61f8349dd5fc6,
64'h1e55b052fdb2e2c5,64'h4bd6bb172e15d48c,64'h6564115e40c74369,64'h0001000000000000,
64'h52a870c4a011519b,64'ha6b394600e9ca35c,64'hc462328a529393c6,64'hb2a043752e8cf9ac,
64'hbf8d789c65167b66,64'hfcb53e480f78671b,64'hd13a7a8ad82139a2,64'hfffffdfefe000201,
64'h98bdc1d5572091a2,64'h77dc1642a8ddef0c,64'h10f99eea89fc23c0,64'h2e30fc204eeafe2a,
64'hf2ad8297ed971628,64'h5eb5d8bb70aea45e,64'h2b208af5063a1b45,64'h0008000000000000,
64'h95438627008a8cd6,64'h359ca30574e51adb,64'h23119458949c9e2a,64'h95021bae7467cd5b,
64'hfc6bc4e828b3db2b,64'he5a9f2477bc338d1,64'h89d3d45cc109cd0a,64'hffffeffef0001001,
64'hc5ee0eaeb9048d0c,64'hbee0b21846ef785d,64'h87ccf7544fe11e00,64'h7187e1037757f14f,
64'h956c14c66cb8b139,64'hf5aec5dd857522ee,64'h590457a931d0da27,64'h0040000000000000,
64'haa1c313c045466ac,64'hace5182ca728d6d7,64'h188ca2c5a4e4f14f,64'ha810dd77a33e6ad4,
64'he35e2748459ed951,64'h2d4f9242de19c681,64'h4e9ea2ea084e684c,64'hffff7ffe80008001,
64'h2f70757bc824685a,64'hf70590c7377bc2e3,64'h3e67baa67f08effc,64'h8c3f081ebabf8a75,
64'hab60a63765c589c4,64'had762ef32ba91769,64'hc822bd4b8e86d136,64'h0200000000000000,
64'h50e189e522a3355b,64'h6728c16a3946b6b3,64'hc465162d27278a78,64'h4086ebc219f3569b,
64'h1af13a492cf6ca81,64'h6a7c9217f0ce3407,64'h74f517524273425e,64'hfffbfffb00040001,
64'h7b83abdf412342cf,64'hb82c8640bbde1711,64'hf33dd534f8477fdf,64'h61f840f9d5fc53a4,
64'h5b0531c02e2c4e1b,64'h6bb1779e5d48bb43,64'h4115ea62743689aa,64'h1000000000000000,
64'h870c4f2b1519aad6,64'h39460b54ca35b595,64'h2328b16f393c53ba,64'h04375e12cf9ab4d6,
64'hd789d24967b65408,64'h53e490c28671a035,64'ha7a8ba95139a12ed,64'hffdfffdf00200001,
64'hdc1d5efd091a1675,64'hc164320adef0b883,64'h99eea9aec23bfef1,64'h0fc207d1afe29d1d,
64'hd8298e03716270d6,64'h5d8bbcf5ea45da15,64'h08af5315a1b44d4e,64'h8000000000000000,
64'h3862795ca8cd56ac,64'hca305aa751adaca7,64'h19458b7ac9e29dcf,64'h21baf0967cd5a6b0,
64'hbc4e92513db2a03a,64'h9f248616338d01a6,64'h3d45d4ad9cd09763,64'hfefffeff01000001,
64'he0eaf7ee48d0b3a2,64'h0b21905cf785c412,64'hcf754d7a11dff784,64'h7e103e8d7f14e8e8,
64'hc14c70218b1386aa,64'hec5de7b1522ed0a6,64'h457a98ad0da26a70,64'h00000003fffffffc,
64'hc313cae6466ab55f,64'h5182d5408d6d6532,64'hca2c5bd64f14ee78,64'h0dd784b4e6ad357f,
64'he274928eed9501cb,64'hf92430b59c680d2c,64'hea2ea56de684bb17,64'hf7fff7ff08000001,
64'h0757bf7946859d09,64'h590c82e7bc2e2090,64'h7baa6bd68effbc1a,64'hf081f46ef8a7473d,
64'h0a638112589c354a,64'h62ef3d9191768529,64'h2bd4c56a6d13537e,64'h0000001fffffffe0,
64'h189e57383355aaf2,64'h8c16aa066b6b298e,64'h5162deb878a773ba,64'h6ebc25a73569abf8,
64'h13a4947e6ca80e51,64'hc92185b3e3406959,64'h51752b763425d8b1,64'hbfffbfff40000001,
64'h3abdfbca342ce848,64'hc864173fe171047e,64'hdd535eb777fde0cd,64'h840fa37ec53a39e1,
64'h531c0892c4e1aa50,64'h1779ec8f8bb42945,64'h5ea62b54689a9bef,64'h000000ffffffff00,
64'hc4f2b9c19aad5790,64'h60b550375b594c6c,64'h8b16f5c5c53b9dce,64'h75e12d3cab4d5fbd,
64'h9d24a3f365407288,64'h490c2da51a034ac2,64'h8ba95bb3a12ec586,64'hfffdffff00000003,
64'hd5efde52a167423f,64'h4320ba050b8823ea,64'hea9af5c1bfef0662,64'h207d1bfa29d1cf04,
64'h98e04498270d527e,64'hbbcf647c5da14a28,64'hf5315aa544d4df76,64'h000007fffffff800,
64'h2795ce12d56abc7a,64'h05aa81bddaca635d,64'h58b7ae3229dcee6c,64'haf0969e85a6afde5,
64'he9251f9f2a03943c,64'h48616d2ad01a560e,64'h5d4adda109762c2c,64'hffefffff00000011,
64'haf7ef29b0b3a11f2,64'h1905d02a5c411f4e,64'h54d7ae14ff783309,64'h03e8dfd24e8e781f,
64'hc70224c5386a93ec,64'hde7b23e7ed0a513b,64'ha98ad53126a6fba9,64'h00003fffffffc000,
64'h3cae7097ab55e3cf,64'h2d540deed6531ae8,64'hc5bd71934ee7735e,64'h784b4f47d357ef23,
64'h4928fd00501ca1d9,64'h430b695880d2b06e,64'hea56ed0a4bb1615e,64'hff7fffff00000081,
64'h7bf794dd59d08f8b,64'hc82e8152e208fa70,64'ha6bd70a9fbc19846,64'h1f46fe927473c0f8,
64'h3811262fc3549f5a,64'hf3d91f45685289d2,64'h4c56a98e3537dd43,64'h0001fffffffe0000,
64'he57384be5aaf1e77,64'h6aa06f77b298d73f,64'h2deb8ca0773b9aea,64'hc25a7a419abf7915,
64'h4947e80480e50ec6,64'h185b4ac60695836e,64'h52b768595d8b0ae9,64'hfbffffff00000401,
64'hdfbca6edce847c55,64'h41740a9d1047d37a,64'h35eb8554de0cc22b,64'hfa37f493a39e07c0,
64'hc089317f1aa4facf,64'h9ec8fa3242944e89,64'h62b54c73a9beea16,64'h000ffffffff00000,
64'h2b9c25f9d578f3b1,64'h55037bc094c6b9f5,64'h6f5c6504b9dcd74f,64'h12d3d212d5fbc8a2,
64'h4a3f40260728762e,64'hc2da563034ac1b70,64'h95bb42ccec585746,64'hdfffffff00002001,
64'hfde537747423e2a2,64'h0ba054ea823e9bce,64'haf5c2aa7f0661157,64'hd1bfa4a41cf03df9,
64'h04498bfed527d672,64'hf647d19614a27444,64'h15aa63a04df750ad,64'h007fffffff800000,
64'h5ce12fcfabc79d87,64'ha81bde06a635cfa6,64'h7ae32828cee6ba75,64'h969e9096afde4510,
64'h51fa01323943b16e,64'h16d2b187a560db7a,64'hadda166b62c2ba2c,64'hfffffffe00010002,
64'hef29bbaaa11f1509,64'h5d02a75411f4de70,64'h7ae1554483308ab3,64'h8dfd2526e781efc2,
64'h224c5ff6a93eb390,64'hb23e8cb7a513a219,64'had531d026fba8568,64'h03fffffffc000000,
64'he7097e7f5e3cec36,64'h40def03a31ae7d2b,64'hd71941497735d3a5,64'hb4f484b97ef2287c,
64'h8fd00993ca1d8b6e,64'hb6958c3d2b06dbd0,64'h6ed0b3601615d15b,64'hfffffff700080009,
64'h794ddd5c08f8a841,64'he8153aa28fa6f37e,64'hd70aaa2719845595,64'h6fe9293b3c0f7e0c,
64'h1262ffb649f59c7f,64'h91f465c2289d10c3,64'h6a98e8187dd42b3b,64'h1fffffffe0000000,
64'h384bf401f1e761a9,64'h06f781d38d73e956,64'hb8ca0a51b9ae9d22,64'ha7a425d0f79143db,
64'h7e804ca250ec5b6c,64'hb4ac61ee5836de7b,64'h76859b03b0ae8ad5,64'hffffffbf00400041,
64'hca6eeae347c54205,64'h40a9d51b7d379be9,64'hb855513ecc22aca2,64'h7f4949dce07bf05d,
64'h9317fdb24face3f8,64'h8fa32e1544e88614,64'h54c740c6eea159d5,64'hffffffff00000000,
64'hc25fa0108f3b0d47,64'h37bc0e9c6b9f4ab0,64'hc6505292cd74e90b,64'h3d212e8cbc8a1ed3,
64'hf40265158762db5d,64'ha5630f77c1b6f3d3,64'hb42cd820857456a5,64'hfffffdff02000201,
64'h537757203e2a1022,64'h054ea8dde9bcdf46,64'hc2aa89fb6115650b,64'hfa4a4eea03df82e5,
64'h98bfed967d671fbc,64'h7d1970ae2744309c,64'ha63a0639750acea6,64'hfffffffefffffff9,
64'h12fd008a79d86a32,64'hbde074e45cfa557f,64'h3282949c6ba74852,64'he9097466e450f697,
64'ha01328b33b16dae1,64'h2b187bc30db79e93,64'ha166c1092ba2b523,64'hffffefff10001001,
64'h9bbab903f150810e,64'h2a7546ef4de6fa30,64'h15544fe108ab2852,64'hd25277571efc1721,
64'hc5ff6cb7eb38fddc,64'he8cb85743a2184dd,64'h31d031d0a856752b,64'hfffffffeffffffc1,
64'h97e80453cec35190,64'hef03a727e7d2abf3,64'h9414a4e45d3a428f,64'h484ba33e2287b4b1,
64'h0099459ed8b6d703,64'h58c3de196dbcf497,64'h0b36084e5d15a913,64'hffff7fff80008001,
64'hddd5c8238a84086c,64'h53aa377b6f37d17f,64'haaa27f0845594290,64'h9293babef7e0b902,
64'h2ffb65c559c7eeda,64'h465c2ba8d10c26e1,64'h8e818e8642b3a957,64'hfffffffefffffe01,
64'hbf4022a2761a8c7c,64'h781d39463e955f91,64'ha0a52726e9d21474,64'h425d19f3143da586,
64'h04ca2cf6c5b6b818,64'hc61ef0cd6de7a4b6,64'h59b04272e8ad4898,64'hfffc000300040001,
64'heeae41225420435a,64'h9d51bbdd79be8bf6,64'h5513f8472aca147b,64'h949dd5fbbf05c80c,
64'h7fdb2e2bce3f76cf,64'h32e15d4888613706,64'h740c7436159d4ab4,64'hfffffffefffff001,
64'hfa011518b0d463db,64'hc0e9ca34f4aafc85,64'h0529393c4e90a39b,64'h12e8cf9aa1ed2c2e,
64'h265167b62db5c0c0,64'h30f786716f3d25aa,64'hcd821399456a44be,64'hffe0001f00200001,
64'h75720919a1021ac9,64'hea8ddeefcdf45fac,64'ha89fc23b5650a3d6,64'ha4eeafe1f82e405c,
64'hfed9716171fbb675,64'h970aea454309b82f,64'ha063a1b3acea559d,64'hfffffffeffff8001,
64'hd008a8cc86a31ed1,64'h074e51ada557e422,64'h2949c9e274851cd8,64'h97467cd50f696170,
64'h328b3db26dae05ff,64'h87bc338c79e92d4f,64'h6c109cd02b5225ea,64'hff0000ff01000001,
64'hab9048d00810d645,64'h546ef7856fa2fd59,64'h44fe11dfb2851eab,64'h27757f14c17202db,
64'hf6cb8b128fddb3a1,64'hb857522e184dc174,64'h031d0da26752ace3,64'hfffffffefffc0001,
64'h8045466a3518f682,64'h3a728d6d2abf2110,64'h4a4e4f14a428e6bf,64'hba33e6ac7b4b0b7c,
64'h9459ed946d702ff7,64'h3de19c67cf496a74,64'h6084e6845a912f4d,64'hf80007ff08000001,
64'h5c8246854086b223,64'ha377bc2d7d17eac6,64'h27f08eff9428f556,64'h3babf8a70b9016d7,
64'hb65c589b7eed9d01,64'hc2ba9175c26e0b9b,64'h18e86d133a956718,64'hfffffffeffe00001,
64'h022a3355a8c7b40c,64'hd3946b6a55f9087f,64'h527278a7214735f6,64'hd19f3568da585bdb,
64'ha2cf6ca76b817fb4,64'hef0ce33f7a4b539f,64'h04273425d4897a65,64'hc0003fff40000001,
64'he412342c04359116,64'h1bbde170e8bf562b,64'h3f8477fda147aaaf,64'hdd5fc5395c80b6b7,
64'hb2e2c4e0f76ce803,64'h15d48bb413705cd2,64'hc7436899d4ab38c0,64'hfffffffeff000001,
64'h11519aad463da060,64'h9ca35b58afc843f2,64'h9393c53b0a39afae,64'h8cf9ab4cd2c2ded2,
64'h167b65405c0bfd9b,64'h78671a02d25a9cf1,64'h2139a12ea44bd328,64'h0002000000000002,
64'h2091a16721ac88a9,64'hddef0b8745fab158,64'hfc23bfee0a3d5577,64'heafe29d0e405b5b2,
64'h9716270cbb674013,64'haea45da09b82e690,64'h3a1b44d4a559c5fa,64'hfffffffef8000001,
64'h8a8cd56a31ed0300,64'he51adac97e421f8c,64'h9c9e29dc51cd7d6c,64'h67cd5a6a9616f68c,
64'hb3db2a02e05fecd8,64'hc338d01992d4e785,64'h09cd0976225e993f,64'h0010000000000010,
64'h048d0b3a0d644547,64'hef785c402fd58aba,64'he11dff7751eaabb1,64'h57f14e8e202dad89,
64'hb8b13869db3a0094,64'h7522ed09dc17347b,64'hd0da26a62ace2fcf,64'hfffffffec0000001,
64'h5466ab558f6817fc,64'h28d6d652f210fc59,64'he4f14ee68e6beb5c,64'h3e6ad357b0b7b45d,
64'h9ed9501c02ff66bb,64'h19c680d296a73c22,64'h4e684bb112f4c9f8,64'h0080000000000080,
64'h246859d06b222a38,64'h7bc2e2087eac55c9,64'h08effbc18f555d81,64'hbf8a7473016d6c46,
64'hc589c353d9d0049b,64'ha9176851e0b9a3d5,64'h86d1353756717e72,64'hfffffffd00000001,
64'ha3355aae7b40bfde,64'h46b6b2989087e2c7,64'h278a773b735f5ad9,64'hf3569abe85bda2e7,
64'hf6ca80e417fb35d4,64'hce340694b539e110,64'h73425d8a97a64fbe,64'h0400000000000400,
64'h2342ce84591151bf,64'hde171046f562ae45,64'h477fde0c7aaaec08,64'hfc53a39d0b6b622b,
64'h2c4e1aa4ce8024d2,64'h48bb429405cd1ea3,64'h3689a9beb38bf38c,64'hffffffef00000001,
64'h19aad578da05feeb,64'h35b594c6843f1636,64'h3c53b9dc9afad6c7,64'h9ab4d5fb2ded1731,
64'hb6540727bfd9ae99,64'h71a034aba9cf087a,64'h9a12ec57bd327ded,64'h2000000000002000,
64'h1a167423c88a8df7,64'hf0b8823dab157222,64'h3bfef065d557603e,64'he29d1cef5b5b1151,
64'h6270d5277401268f,64'h45da14a22e68f516,64'hb44d4df69c5f9c5f,64'hffffff7f00000001,
64'hcd56abc6d02ff758,64'hadaca63521f8b1af,64'he29dcee5d7d6b637,64'hd5a6afdd6f68b984,
64'hb2a03942fecd74c3,64'h8d01a5604e7843cd,64'hd09762c1e993ef64,64'h000000010000ffff,
64'hd0b3a11e44546fb8,64'h85c411f458ab9109,64'hdff7832faabb01ef,64'h14e8e781dad88a81,
64'h1386a93ea0093475,64'h2ed0a5137347a8ae,64'ha26a6fb9e2fce2f3,64'hfffffbff00000001,
64'h6ab55e3c817fbaba,64'h6d6531ae0fc58d73,64'h14ee7735beb5b1b1,64'had357ef17b45cc1a,
64'h9501ca1cf66ba613,64'h680d2b0673c21e64,64'h84bb16154c9f7b1a,64'h000000080007fff8,
64'h859d08f822a37dba,64'h2e208fa6c55c8844,64'hffbc198355d80f72,64'ha7473c0ed6c45408,
64'h9c3549f50049a3a8,64'h7685289c9a3d456f,64'h13537dd417e71793,64'hffffdfff00000001,
64'h55aaf1e70bfdd5cd,64'h6b298d737e2c6b95,64'ha773b9adf5ad8d88,64'h69abf790da2e60cb,
64'ha80e50ebb35d3094,64'h406958369e10f31d,64'h25d8b0ae64fbd8cc,64'h00000040003fffc0,
64'h2ce847c5151bedcc,64'h71047d372ae4421f,64'hfde0cc21aec07b89,64'h3a39e07bb622a03b,
64'he1aa4fac024d1d3c,64'hb42944e7d1ea2b75,64'h9a9beea0bf38bc98,64'hfffeffff00000001,
64'had578f3a5feeae66,64'h594c6b9ef1635ca5,64'h3b9dcd74ad6c6c3b,64'h4d5fbc89d1730655,
64'h407287629ae9849b,64'h034ac1b6f08798e6,64'h2ec5857427dec65f,64'h0000020001fffe00,
64'h67423e29a8df6e5f,64'h8823e9bc572210f5,64'hef0661147603dc41,64'hd1cf03deb11501d7,
64'h0d527d671268e9d9,64'ha14a27438f515ba3,64'hd4df7509f9c5e4bc,64'hfff7ffff00000001,
64'h6abc79d7ff75732b,64'hca635cf98b1ae526,64'hdcee6ba66b6361d7,64'h6afde4508b9832a6,
64'h03943b16d74c24d6,64'h1a560db7843cc730,64'h762c2ba23ef632f7,64'h000010000ffff000,
64'h3a11f15046fb72f5,64'h411f4de6b91087a4,64'h783308aab01ee201,64'h8e781efb88a80eb2,
64'h6a93eb3893474ec8,64'h0a513a217a8add13,64'ha6fba855ce2f25da,64'hffbfffff00000001,
64'h55e3cec2fbab9955,64'h531ae7d258d7292a,64'he7735d395b1b0eb2,64'h57ef22875cc1952d,
64'h1ca1d8b6ba6126b0,64'hd2b06dbc21e63980,64'hb1615d14f7b197b5,64'h000080007fff8000,
64'hd08f8a8337db97a7,64'h08fa6f37c8843d1e,64'hc198455880f71005,64'h73c0f7e04540758c,
64'h549f59c79a3a763d,64'h5289d10bd456e898,64'h37dd42b371792ecb,64'hfdffffff00000001,
64'haf1e7619dd5ccaa6,64'h98d73e94c6b9494e,64'h3b9ae9d1d8d87589,64'hbf79143ce60ca966,
64'he50ec5b5d3093580,64'h95836de70f31cbfa,64'h8b0ae8acbd8cbda3,64'h00040003fffc0000,
64'h847c541fbedcbd32,64'h47d379be4421e8f0,64'h0cc22aca07b88022,64'h9e07bf052a03ac5d,
64'ha4face3ed1d3b1e6,64'h944e8860a2b744be,64'hbeea159c8bc97657,64'hefffffff00000001,
64'h78f3b0d3eae6552b,64'hc6b9f4aa35ca4a6c,64'hdcd74e8fc6c3ac47,64'hfbc8a1ec30654b2b,
64'h28762db59849abf9,64'hac1b6f3c798e5fcc,64'h58574569ec65ed14,64'h0020001fffe00000,
64'h23e2a101f6e5e98c,64'h3e9bcdf4210f477e,64'h661156503dc40110,64'hf03df82d501d62e4,
64'h27d671fb8e9d8f2b,64'ha274430915ba25ec,64'hf750ace95e4bb2b3,64'h7fffffff00000001,
64'hc79d86a25732a955,64'h35cfa557ae52535a,64'he6ba7484361d6232,64'hde450f68832a5951,
64'h43b16dadc24d5fc7,64'h60db79e8cc72fe5b,64'hc2ba2b51632f689e,64'h010000ffff000000,
64'h1f150810b72f4c5f,64'hf4de6fa2087a3bef,64'h308ab284ee20087d,64'h81efc17180eb1719,
64'h3eb38fdd74ec7957,64'h13a2184dadd12f5b,64'hba856751f25d9591,64'hfffffffb00000005,
64'h3cec3518b9954aa2,64'hae7d2abe72929acf,64'h35d3a428b0eb1189,64'hf2287b4a1952ca82,
64'h1d8b6d70126afe36,64'h06dbcf496397f2d5,64'h15d15a91197b44ea,64'h080007fff8000000,
64'hf8a84085b97a62f8,64'ha6f37d1743d1df71,64'h84559428710043e7,64'h0f7e0b900758b8c4,
64'hf59c7eeca763cab7,64'h9d10c26d6e897ad8,64'hd42b3a9492ecac83,64'hffffffdf00000021,
64'he761a8c6ccaa550f,64'h73e955f89494d673,64'hae9d214687588c47,64'h9143da57ca965409,
64'hec5b6b809357f1b0,64'h36de7a4b1cbf96a8,64'hae8ad488cbda2750,64'h40003fffc0000000,
64'hc5420434cbd317b9,64'h379be8bf1e8efb83,64'h22aca14788021f34,64'h7bf05c803ac5c620,
64'hace3f76c3b1e55b1,64'he886136f744bd6bc,64'ha159d4aa97656412,64'hfffffeff00000101,
64'h3b0d463d6552a871,64'h9f4aafc7a4a6b395,64'h74e90a393ac46233,64'h8a1ed2c254b2a044,
64'h62db5c0b9abf8d79,64'hb6f3d259e5fcb53f,64'h7456a44b5ed13a7b,64'h0001fffffffffffe,
64'h2a1021ac5e98bdc2,64'hbcdf45f9f477dc17,64'h15650a3d4010f99f,64'hdf82e404d62e30fd,
64'h671fbb66d8f2ad83,64'h44309b82a25eb5d9,64'h0acea559bb2b208b,64'hfffff7ff00000801,
64'hd86a31ec2a954387,64'hfa557e4125359ca4,64'ha74851ccd6231195,64'h50f69616a595021c,
64'h16dae05fd5fc6bc5,64'hb79e92d42fe5a9f3,64'ha2b5225df689d3d5,64'h000ffffffffffff0,
64'h50810d63f4c5ee0f,64'he6fa2fd4a3bee0b3,64'hab2851ea0087ccf8,64'hfc17202cb17187e2,
64'h38fddb39c7956c15,64'h2184dc1712f5aec6,64'h56752acdd9590458,64'hffffbfff00004001,
64'hc3518f6754aa1c32,64'hd2abf21029ace519,64'h3a428e6bb1188ca3,64'h87b4b0b72ca810de,
64'hb6d702feafe35e28,64'hbcf496a67f2d4f93,64'h15a912f4b44e9ea3,64'h007fffffffffff80,
64'h84086b21a62f7076,64'h37d17eac1df70591,64'h59428f55043e67bb,64'he0b9016c8b8c3f09,
64'hc7eed9cf3cab60a7,64'h0c26e0b997ad762f,64'hb3a95670cac822be,64'hfffdffff00020001,
64'h1a8c7b40a550e18a,64'h955f90874d6728c2,64'hd214735e88c46517,64'h3da585bd654086ec,
64'hb6b817fa7f1af13b,64'he7a4b538f96a7c93,64'had4897a5a274f518,64'h03fffffffffffc00,
64'h20435911317b83ac,64'hbe8bf561efb82c87,64'hca147aaa21f33dd6,64'h05c80b6b5c61f841,
64'h3f76ce7fe55b0532,64'h613705ccbd6bb178,64'h9d4ab38b564115eb,64'hffefffff00100001,
64'hd463da052a870c50,64'haafc843e6b39460c,64'h90a39afa462328b2,64'hed2c2dec2a04375f,
64'hb5c0bfd8f8d789d3,64'h3d25a9cecb53e491,64'h6a44bd3213a7a8bb,64'h1fffffffffffe000,
64'h021ac88a8bdc1d5f,64'hf45fab147dc16433,64'h50a3d5570f99eeaa,64'h2e405b5ae30fc208,
64'hfbb674002ad8298f,64'h09b82e68eb5d8bbd,64'hea559c5eb208af54,64'hff7fffff00800001,
64'ha31ed02f5438627a,64'h57e421f859ca305b,64'h851cd7d63119458c,64'h69616f685021baf1,
64'hae05feccc6bc4e93,64'he92d4e775a9f2487,64'h5225e9939d3d45d5,64'h00000000fffeffff,
64'h10d644545ee0eaf8,64'ha2fd58aaee0b2191,64'h851eaaba7ccf754e,64'h7202dad8187e103f,
64'hddb3a00856c14c71,64'h4dc173475aec5de8,64'h52ace2fc90457a99,64'hfbffffff04000001,
64'h18f6817fa1c313cb,64'hbf210fc4ce5182d6,64'h28e6beb588ca2c5c,64'h4b0b7b45810dd785,
64'h702ff66b35e27493,64'h496a73c1d4f92431,64'h912f4c9ee9ea2ea6,64'h00000007fff7fff8,
64'h86b222a2f70757c0,64'h17eac55c70590c83,64'h28f555d7e67baa6c,64'h9016d6c3c3f081f5,
64'hed9d0048b60a6382,64'h6e0b9a3cd762ef3e,64'h956717e6822bd4c6,64'hdfffffff20000001,
64'hc7b40bfd0e189e58,64'hf9087e2b728c16ab,64'h4735f5ad465162df,64'h585bda2e086ebc26,
64'h817fb35caf13a495,64'h4b539e10a7c92186,64'h897a64fb4f51752c,64'h0000003fffbfffc0,
64'h3591151bb83abdfc,64'hbf562ae382c86418,64'h47aaaec033dd535f,64'h80b6b6221f840fa4,
64'h6ce8024cb0531c09,64'h705cd1e9bb1779ed,64'hab38bf38115ea62c,64'h0000000000000001
};
  //------------------------
  // 256
  //------------------------
  localparam [2*256-1:0][63:0] NTT_GF64_BWD_N256_PHI_L = {
64'hc843f1629460b551,64'hc2ded1724375e12e,64'h5a9cf0873e490c2e,64'h000001fffdfffe00,
64'hfab15721164320bb,64'h05b5b114fc207d1c,64'h82e68f50d8bbcf65,64'h0000000000000008,
64'h421f8b1aa305aa82,64'h16f68b981baf096a,64'hd4e7843bf248616e,64'h00000fffeffff000,
64'hd58ab90fb21905d1,64'h2dad88a7e103e8e0,64'h17347a8ac5de7b24,64'h0000000000000040,
64'h10fc58d7182d540e,64'hb7b45cc0dd784b50,64'ha73c21e592430b6a,64'h00007fff7fff8000,
64'hac55c88390c82e82,64'h6d6c4540081f46ff,64'hb9a3d4562ef3d920,64'h0000000000000200,
64'h87e2c6b8c16aa070,64'hbda2e60bebc25a7b,64'h39e10f3192185b4b,64'h0003fffbfffc0000,
64'h62ae44218641740b,64'h6b622a0340fa37f5,64'hcd1ea2b6779ec8fb,64'h0000000000001000,
64'h3f1635ca0b55037c,64'hed1730645e12d3d3,64'hcf08798d90c2da57,64'h001fffdfffe00000,
64'h1572210f320ba055,64'h5b11501d07d1bfa5,64'h68f515b9bcf647d2,64'h0000000000008000,
64'hf8b1ae515aa81bdf,64'h68b98329f0969e91,64'h7843cc728616d2b2,64'h00fffeffff000000,
64'hab910879905d02a8,64'hd88a80ea3e8dfd26,64'h47a8add0e7b23e8d,64'h0000000000040000,
64'hc58d7291d540def1,64'h45cc195284b4f485,64'hc21e639730b6958d,64'h07fff7fff8000000,
64'h5c8843d182e8153b,64'hc4540757f46fe92a,64'h3d456e893d91f466,64'h0000000000200000,
64'h2c6b9494aa06f782,64'h2e60ca9625a7a426,64'h10f31cbf85b4ac62,64'h3fffbfffc0000000,
64'he4421e8e1740a9d6,64'h22a03ac5a37f494a,64'hea2b744aec8fa32f,64'h0000000001000000,
64'h635ca4a65037bc0f,64'h730654b22d3d212f,64'h8798e5fc2da56310,64'hfffdfffeffffffff,
64'h2210f477ba054ea9,64'h1501d62e1bfa4a4f,64'h515ba25e647d1971,64'h0000000008000000,
64'h1ae5253581bde075,64'h9832a59469e90975,64'h3cc72fe56d2b187c,64'hffeffffefffffff1,
64'h1087a3bed02a7547,64'ha80eb170dfd25278,64'h8add12f523e8cb86,64'h0000000040000000,
64'hd72929ac0def03a8,64'hc1952ca74f484ba4,64'he6397f2c6958c3df,64'hff7ffffeffffff81,
64'h843d1df68153aa38,64'h40758b8bfe9293bb,64'h56e897ad1f465c2c,64'h0000000200000000,
64'hb9494d666f781d3a,64'h0ca965407a425d1a,64'h31cbf96a4ac61ef1,64'hfbfffffefffffc01,
64'h21e8efb80a9d51bc,64'h03ac5c61f4949dd6,64'hb744bd6afa32e15e,64'h0000001000000000,
64'hca4a6b387bc0e9cb,64'h654b2a03d212e8d0,64'h8e5fcb535630f787,64'hdffffffeffffe001,
64'h0f477dc154ea8ddf,64'h1d62e30fa4a4eeb0,64'hba25eb5cd1970aeb,64'h0000008000000000,
64'h525359c9de074e52,64'h2a5950219097467d,64'h72fe5a9eb187bc34,64'hfffffffdffff0002,
64'h7a3bee0aa7546ef8,64'heb17187d25277580,64'hd12f5aeb8cb85753,64'h0000040000000000,
64'h929ace50f03a728e,64'h52ca810d84ba33e7,64'h97f2d4f88c3de19d,64'hfffffff6fff80009,
64'hd1df70583aa377bd,64'h58b8c3f0293babf9,64'h897ad76265c2ba92,64'h0000200000000000,
64'h94d6728b81d3946c,64'h9654086e25d19f36,64'hbf96a7c861ef0ce4,64'hffffffbeffc00041,
64'h8efb82c7d51bbde2,64'hc5c61f8349dd5fc6,64'h4bd6bb172e15d48c,64'h0001000000000000,
64'ha6b394600e9ca35c,64'hb2a043752e8cf9ac,64'hfcb53e480f78671b,64'hfffffdfefe000201,
64'h77dc1642a8ddef0c,64'h2e30fc204eeafe2a,64'h5eb5d8bb70aea45e,64'h0008000000000000,
64'h359ca30574e51adb,64'h95021bae7467cd5b,64'he5a9f2477bc338d1,64'hffffeffef0001001,
64'hbee0b21846ef785d,64'h7187e1037757f14f,64'hf5aec5dd857522ee,64'h0040000000000000,
64'hace5182ca728d6d7,64'ha810dd77a33e6ad4,64'h2d4f9242de19c681,64'hffff7ffe80008001,
64'hf70590c7377bc2e3,64'h8c3f081ebabf8a75,64'had762ef32ba91769,64'h0200000000000000,
64'h6728c16a3946b6b3,64'h4086ebc219f3569b,64'h6a7c9217f0ce3407,64'hfffbfffb00040001,
64'hb82c8640bbde1711,64'h61f840f9d5fc53a4,64'h6bb1779e5d48bb43,64'h1000000000000000,
64'h39460b54ca35b595,64'h04375e12cf9ab4d6,64'h53e490c28671a035,64'hffdfffdf00200001,
64'hc164320adef0b883,64'h0fc207d1afe29d1d,64'h5d8bbcf5ea45da15,64'h8000000000000000,
64'hca305aa751adaca7,64'h21baf0967cd5a6b0,64'h9f248616338d01a6,64'hfefffeff01000001,
64'h0b21905cf785c412,64'h7e103e8d7f14e8e8,64'hec5de7b1522ed0a6,64'h00000003fffffffc,
64'h5182d5408d6d6532,64'h0dd784b4e6ad357f,64'hf92430b59c680d2c,64'hf7fff7ff08000001,
64'h590c82e7bc2e2090,64'hf081f46ef8a7473d,64'h62ef3d9191768529,64'h0000001fffffffe0,
64'h8c16aa066b6b298e,64'h6ebc25a73569abf8,64'hc92185b3e3406959,64'hbfffbfff40000001,
64'hc864173fe171047e,64'h840fa37ec53a39e1,64'h1779ec8f8bb42945,64'h000000ffffffff00,
64'h60b550375b594c6c,64'h75e12d3cab4d5fbd,64'h490c2da51a034ac2,64'hfffdffff00000003,
64'h4320ba050b8823ea,64'h207d1bfa29d1cf04,64'hbbcf647c5da14a28,64'h000007fffffff800,
64'h05aa81bddaca635d,64'haf0969e85a6afde5,64'h48616d2ad01a560e,64'hffefffff00000011,
64'h1905d02a5c411f4e,64'h03e8dfd24e8e781f,64'hde7b23e7ed0a513b,64'h00003fffffffc000,
64'h2d540deed6531ae8,64'h784b4f47d357ef23,64'h430b695880d2b06e,64'hff7fffff00000081,
64'hc82e8152e208fa70,64'h1f46fe927473c0f8,64'hf3d91f45685289d2,64'h0001fffffffe0000,
64'h6aa06f77b298d73f,64'hc25a7a419abf7915,64'h185b4ac60695836e,64'hfbffffff00000401,
64'h41740a9d1047d37a,64'hfa37f493a39e07c0,64'h9ec8fa3242944e89,64'h000ffffffff00000,
64'h55037bc094c6b9f5,64'h12d3d212d5fbc8a2,64'hc2da563034ac1b70,64'hdfffffff00002001,
64'h0ba054ea823e9bce,64'hd1bfa4a41cf03df9,64'hf647d19614a27444,64'h007fffffff800000,
64'ha81bde06a635cfa6,64'h969e9096afde4510,64'h16d2b187a560db7a,64'hfffffffe00010002,
64'h5d02a75411f4de70,64'h8dfd2526e781efc2,64'hb23e8cb7a513a219,64'h03fffffffc000000,
64'h40def03a31ae7d2b,64'hb4f484b97ef2287c,64'hb6958c3d2b06dbd0,64'hfffffff700080009,
64'he8153aa28fa6f37e,64'h6fe9293b3c0f7e0c,64'h91f465c2289d10c3,64'h1fffffffe0000000,
64'h06f781d38d73e956,64'ha7a425d0f79143db,64'hb4ac61ee5836de7b,64'hffffffbf00400041,
64'h40a9d51b7d379be9,64'h7f4949dce07bf05d,64'h8fa32e1544e88614,64'hffffffff00000000,
64'h37bc0e9c6b9f4ab0,64'h3d212e8cbc8a1ed3,64'ha5630f77c1b6f3d3,64'hfffffdff02000201,
64'h054ea8dde9bcdf46,64'hfa4a4eea03df82e5,64'h7d1970ae2744309c,64'hfffffffefffffff9,
64'hbde074e45cfa557f,64'he9097466e450f697,64'h2b187bc30db79e93,64'hffffefff10001001,
64'h2a7546ef4de6fa30,64'hd25277571efc1721,64'he8cb85743a2184dd,64'hfffffffeffffffc1,
64'hef03a727e7d2abf3,64'h484ba33e2287b4b1,64'h58c3de196dbcf497,64'hffff7fff80008001,
64'h53aa377b6f37d17f,64'h9293babef7e0b902,64'h465c2ba8d10c26e1,64'hfffffffefffffe01,
64'h781d39463e955f91,64'h425d19f3143da586,64'hc61ef0cd6de7a4b6,64'hfffc000300040001,
64'h9d51bbdd79be8bf6,64'h949dd5fbbf05c80c,64'h32e15d4888613706,64'hfffffffefffff001,
64'hc0e9ca34f4aafc85,64'h12e8cf9aa1ed2c2e,64'h30f786716f3d25aa,64'hffe0001f00200001,
64'hea8ddeefcdf45fac,64'ha4eeafe1f82e405c,64'h970aea454309b82f,64'hfffffffeffff8001,
64'h074e51ada557e422,64'h97467cd50f696170,64'h87bc338c79e92d4f,64'hff0000ff01000001,
64'h546ef7856fa2fd59,64'h27757f14c17202db,64'hb857522e184dc174,64'hfffffffefffc0001,
64'h3a728d6d2abf2110,64'hba33e6ac7b4b0b7c,64'h3de19c67cf496a74,64'hf80007ff08000001,
64'ha377bc2d7d17eac6,64'h3babf8a70b9016d7,64'hc2ba9175c26e0b9b,64'hfffffffeffe00001,
64'hd3946b6a55f9087f,64'hd19f3568da585bdb,64'hef0ce33f7a4b539f,64'hc0003fff40000001,
64'h1bbde170e8bf562b,64'hdd5fc5395c80b6b7,64'h15d48bb413705cd2,64'hfffffffeff000001,
64'h9ca35b58afc843f2,64'h8cf9ab4cd2c2ded2,64'h78671a02d25a9cf1,64'h0002000000000002,
64'hddef0b8745fab158,64'heafe29d0e405b5b2,64'haea45da09b82e690,64'hfffffffef8000001,
64'he51adac97e421f8c,64'h67cd5a6a9616f68c,64'hc338d01992d4e785,64'h0010000000000010,
64'hef785c402fd58aba,64'h57f14e8e202dad89,64'h7522ed09dc17347b,64'hfffffffec0000001,
64'h28d6d652f210fc59,64'h3e6ad357b0b7b45d,64'h19c680d296a73c22,64'h0080000000000080,
64'h7bc2e2087eac55c9,64'hbf8a7473016d6c46,64'ha9176851e0b9a3d5,64'hfffffffd00000001,
64'h46b6b2989087e2c7,64'hf3569abe85bda2e7,64'hce340694b539e110,64'h0400000000000400,
64'hde171046f562ae45,64'hfc53a39d0b6b622b,64'h48bb429405cd1ea3,64'hffffffef00000001,
64'h35b594c6843f1636,64'h9ab4d5fb2ded1731,64'h71a034aba9cf087a,64'h2000000000002000,
64'hf0b8823dab157222,64'he29d1cef5b5b1151,64'h45da14a22e68f516,64'hffffff7f00000001,
64'hadaca63521f8b1af,64'hd5a6afdd6f68b984,64'h8d01a5604e7843cd,64'h000000010000ffff,
64'h85c411f458ab9109,64'h14e8e781dad88a81,64'h2ed0a5137347a8ae,64'hfffffbff00000001,
64'h6d6531ae0fc58d73,64'had357ef17b45cc1a,64'h680d2b0673c21e64,64'h000000080007fff8,
64'h2e208fa6c55c8844,64'ha7473c0ed6c45408,64'h7685289c9a3d456f,64'hffffdfff00000001,
64'h6b298d737e2c6b95,64'h69abf790da2e60cb,64'h406958369e10f31d,64'h00000040003fffc0,
64'h71047d372ae4421f,64'h3a39e07bb622a03b,64'hb42944e7d1ea2b75,64'hfffeffff00000001,
64'h594c6b9ef1635ca5,64'h4d5fbc89d1730655,64'h034ac1b6f08798e6,64'h0000020001fffe00,
64'h8823e9bc572210f5,64'hd1cf03deb11501d7,64'ha14a27438f515ba3,64'hfff7ffff00000001,
64'hca635cf98b1ae526,64'h6afde4508b9832a6,64'h1a560db7843cc730,64'h000010000ffff000,
64'h411f4de6b91087a4,64'h8e781efb88a80eb2,64'h0a513a217a8add13,64'hffbfffff00000001,
64'h531ae7d258d7292a,64'h57ef22875cc1952d,64'hd2b06dbc21e63980,64'h000080007fff8000,
64'h08fa6f37c8843d1e,64'h73c0f7e04540758c,64'h5289d10bd456e898,64'hfdffffff00000001,
64'h98d73e94c6b9494e,64'hbf79143ce60ca966,64'h95836de70f31cbfa,64'h00040003fffc0000,
64'h47d379be4421e8f0,64'h9e07bf052a03ac5d,64'h944e8860a2b744be,64'hefffffff00000001,
64'hc6b9f4aa35ca4a6c,64'hfbc8a1ec30654b2b,64'hac1b6f3c798e5fcc,64'h0020001fffe00000,
64'h3e9bcdf4210f477e,64'hf03df82d501d62e4,64'ha274430915ba25ec,64'h7fffffff00000001,
64'h35cfa557ae52535a,64'hde450f68832a5951,64'h60db79e8cc72fe5b,64'h010000ffff000000,
64'hf4de6fa2087a3bef,64'h81efc17180eb1719,64'h13a2184dadd12f5b,64'hfffffffb00000005,
64'hae7d2abe72929acf,64'hf2287b4a1952ca82,64'h06dbcf496397f2d5,64'h080007fff8000000,
64'ha6f37d1743d1df71,64'h0f7e0b900758b8c4,64'h9d10c26d6e897ad8,64'hffffffdf00000021,
64'h73e955f89494d673,64'h9143da57ca965409,64'h36de7a4b1cbf96a8,64'h40003fffc0000000,
64'h379be8bf1e8efb83,64'h7bf05c803ac5c620,64'he886136f744bd6bc,64'hfffffeff00000101,
64'h9f4aafc7a4a6b395,64'h8a1ed2c254b2a044,64'hb6f3d259e5fcb53f,64'h0001fffffffffffe,
64'hbcdf45f9f477dc17,64'hdf82e404d62e30fd,64'h44309b82a25eb5d9,64'hfffff7ff00000801,
64'hfa557e4125359ca4,64'h50f69616a595021c,64'hb79e92d42fe5a9f3,64'h000ffffffffffff0,
64'he6fa2fd4a3bee0b3,64'hfc17202cb17187e2,64'h2184dc1712f5aec6,64'hffffbfff00004001,
64'hd2abf21029ace519,64'h87b4b0b72ca810de,64'hbcf496a67f2d4f93,64'h007fffffffffff80,
64'h37d17eac1df70591,64'he0b9016c8b8c3f09,64'h0c26e0b997ad762f,64'hfffdffff00020001,
64'h955f90874d6728c2,64'h3da585bd654086ec,64'he7a4b538f96a7c93,64'h03fffffffffffc00,
64'hbe8bf561efb82c87,64'h05c80b6b5c61f841,64'h613705ccbd6bb178,64'hffefffff00100001,
64'haafc843e6b39460c,64'hed2c2dec2a04375f,64'h3d25a9cecb53e491,64'h1fffffffffffe000,
64'hf45fab147dc16433,64'h2e405b5ae30fc208,64'h09b82e68eb5d8bbd,64'hff7fffff00800001,
64'h57e421f859ca305b,64'h69616f685021baf1,64'he92d4e775a9f2487,64'h00000000fffeffff,
64'ha2fd58aaee0b2191,64'h7202dad8187e103f,64'h4dc173475aec5de8,64'hfbffffff04000001,
64'hbf210fc4ce5182d6,64'h4b0b7b45810dd785,64'h496a73c1d4f92431,64'h00000007fff7fff8,
64'h17eac55c70590c83,64'h9016d6c3c3f081f5,64'h6e0b9a3cd762ef3e,64'hdfffffff20000001,
64'hf9087e2b728c16ab,64'h585bda2e086ebc26,64'h4b539e10a7c92186,64'h0000003fffbfffc0,
64'hbf562ae382c86418,64'h80b6b6221f840fa4,64'h705cd1e9bb1779ed,64'h0000000000000001
};
  //------------------------
  // 128
  //------------------------
  localparam [2*128-1:0][63:0] NTT_GF64_BWD_N128_PHI_L = {
64'hc2ded1724375e12e,64'h000001fffdfffe00,64'h05b5b114fc207d1c,64'h0000000000000008,
64'h16f68b981baf096a,64'h00000fffeffff000,64'h2dad88a7e103e8e0,64'h0000000000000040,
64'hb7b45cc0dd784b50,64'h00007fff7fff8000,64'h6d6c4540081f46ff,64'h0000000000000200,
64'hbda2e60bebc25a7b,64'h0003fffbfffc0000,64'h6b622a0340fa37f5,64'h0000000000001000,
64'hed1730645e12d3d3,64'h001fffdfffe00000,64'h5b11501d07d1bfa5,64'h0000000000008000,
64'h68b98329f0969e91,64'h00fffeffff000000,64'hd88a80ea3e8dfd26,64'h0000000000040000,
64'h45cc195284b4f485,64'h07fff7fff8000000,64'hc4540757f46fe92a,64'h0000000000200000,
64'h2e60ca9625a7a426,64'h3fffbfffc0000000,64'h22a03ac5a37f494a,64'h0000000001000000,
64'h730654b22d3d212f,64'hfffdfffeffffffff,64'h1501d62e1bfa4a4f,64'h0000000008000000,
64'h9832a59469e90975,64'hffeffffefffffff1,64'ha80eb170dfd25278,64'h0000000040000000,
64'hc1952ca74f484ba4,64'hff7ffffeffffff81,64'h40758b8bfe9293bb,64'h0000000200000000,
64'h0ca965407a425d1a,64'hfbfffffefffffc01,64'h03ac5c61f4949dd6,64'h0000001000000000,
64'h654b2a03d212e8d0,64'hdffffffeffffe001,64'h1d62e30fa4a4eeb0,64'h0000008000000000,
64'h2a5950219097467d,64'hfffffffdffff0002,64'heb17187d25277580,64'h0000040000000000,
64'h52ca810d84ba33e7,64'hfffffff6fff80009,64'h58b8c3f0293babf9,64'h0000200000000000,
64'h9654086e25d19f36,64'hffffffbeffc00041,64'hc5c61f8349dd5fc6,64'h0001000000000000,
64'hb2a043752e8cf9ac,64'hfffffdfefe000201,64'h2e30fc204eeafe2a,64'h0008000000000000,
64'h95021bae7467cd5b,64'hffffeffef0001001,64'h7187e1037757f14f,64'h0040000000000000,
64'ha810dd77a33e6ad4,64'hffff7ffe80008001,64'h8c3f081ebabf8a75,64'h0200000000000000,
64'h4086ebc219f3569b,64'hfffbfffb00040001,64'h61f840f9d5fc53a4,64'h1000000000000000,
64'h04375e12cf9ab4d6,64'hffdfffdf00200001,64'h0fc207d1afe29d1d,64'h8000000000000000,
64'h21baf0967cd5a6b0,64'hfefffeff01000001,64'h7e103e8d7f14e8e8,64'h00000003fffffffc,
64'h0dd784b4e6ad357f,64'hf7fff7ff08000001,64'hf081f46ef8a7473d,64'h0000001fffffffe0,
64'h6ebc25a73569abf8,64'hbfffbfff40000001,64'h840fa37ec53a39e1,64'h000000ffffffff00,
64'h75e12d3cab4d5fbd,64'hfffdffff00000003,64'h207d1bfa29d1cf04,64'h000007fffffff800,
64'haf0969e85a6afde5,64'hffefffff00000011,64'h03e8dfd24e8e781f,64'h00003fffffffc000,
64'h784b4f47d357ef23,64'hff7fffff00000081,64'h1f46fe927473c0f8,64'h0001fffffffe0000,
64'hc25a7a419abf7915,64'hfbffffff00000401,64'hfa37f493a39e07c0,64'h000ffffffff00000,
64'h12d3d212d5fbc8a2,64'hdfffffff00002001,64'hd1bfa4a41cf03df9,64'h007fffffff800000,
64'h969e9096afde4510,64'hfffffffe00010002,64'h8dfd2526e781efc2,64'h03fffffffc000000,
64'hb4f484b97ef2287c,64'hfffffff700080009,64'h6fe9293b3c0f7e0c,64'h1fffffffe0000000,
64'ha7a425d0f79143db,64'hffffffbf00400041,64'h7f4949dce07bf05d,64'hffffffff00000000,
64'h3d212e8cbc8a1ed3,64'hfffffdff02000201,64'hfa4a4eea03df82e5,64'hfffffffefffffff9,
64'he9097466e450f697,64'hffffefff10001001,64'hd25277571efc1721,64'hfffffffeffffffc1,
64'h484ba33e2287b4b1,64'hffff7fff80008001,64'h9293babef7e0b902,64'hfffffffefffffe01,
64'h425d19f3143da586,64'hfffc000300040001,64'h949dd5fbbf05c80c,64'hfffffffefffff001,
64'h12e8cf9aa1ed2c2e,64'hffe0001f00200001,64'ha4eeafe1f82e405c,64'hfffffffeffff8001,
64'h97467cd50f696170,64'hff0000ff01000001,64'h27757f14c17202db,64'hfffffffefffc0001,
64'hba33e6ac7b4b0b7c,64'hf80007ff08000001,64'h3babf8a70b9016d7,64'hfffffffeffe00001,
64'hd19f3568da585bdb,64'hc0003fff40000001,64'hdd5fc5395c80b6b7,64'hfffffffeff000001,
64'h8cf9ab4cd2c2ded2,64'h0002000000000002,64'heafe29d0e405b5b2,64'hfffffffef8000001,
64'h67cd5a6a9616f68c,64'h0010000000000010,64'h57f14e8e202dad89,64'hfffffffec0000001,
64'h3e6ad357b0b7b45d,64'h0080000000000080,64'hbf8a7473016d6c46,64'hfffffffd00000001,
64'hf3569abe85bda2e7,64'h0400000000000400,64'hfc53a39d0b6b622b,64'hffffffef00000001,
64'h9ab4d5fb2ded1731,64'h2000000000002000,64'he29d1cef5b5b1151,64'hffffff7f00000001,
64'hd5a6afdd6f68b984,64'h000000010000ffff,64'h14e8e781dad88a81,64'hfffffbff00000001,
64'had357ef17b45cc1a,64'h000000080007fff8,64'ha7473c0ed6c45408,64'hffffdfff00000001,
64'h69abf790da2e60cb,64'h00000040003fffc0,64'h3a39e07bb622a03b,64'hfffeffff00000001,
64'h4d5fbc89d1730655,64'h0000020001fffe00,64'hd1cf03deb11501d7,64'hfff7ffff00000001,
64'h6afde4508b9832a6,64'h000010000ffff000,64'h8e781efb88a80eb2,64'hffbfffff00000001,
64'h57ef22875cc1952d,64'h000080007fff8000,64'h73c0f7e04540758c,64'hfdffffff00000001,
64'hbf79143ce60ca966,64'h00040003fffc0000,64'h9e07bf052a03ac5d,64'hefffffff00000001,
64'hfbc8a1ec30654b2b,64'h0020001fffe00000,64'hf03df82d501d62e4,64'h7fffffff00000001,
64'hde450f68832a5951,64'h010000ffff000000,64'h81efc17180eb1719,64'hfffffffb00000005,
64'hf2287b4a1952ca82,64'h080007fff8000000,64'h0f7e0b900758b8c4,64'hffffffdf00000021,
64'h9143da57ca965409,64'h40003fffc0000000,64'h7bf05c803ac5c620,64'hfffffeff00000101,
64'h8a1ed2c254b2a044,64'h0001fffffffffffe,64'hdf82e404d62e30fd,64'hfffff7ff00000801,
64'h50f69616a595021c,64'h000ffffffffffff0,64'hfc17202cb17187e2,64'hffffbfff00004001,
64'h87b4b0b72ca810de,64'h007fffffffffff80,64'he0b9016c8b8c3f09,64'hfffdffff00020001,
64'h3da585bd654086ec,64'h03fffffffffffc00,64'h05c80b6b5c61f841,64'hffefffff00100001,
64'hed2c2dec2a04375f,64'h1fffffffffffe000,64'h2e405b5ae30fc208,64'hff7fffff00800001,
64'h69616f685021baf1,64'h00000000fffeffff,64'h7202dad8187e103f,64'hfbffffff04000001,
64'h4b0b7b45810dd785,64'h00000007fff7fff8,64'h9016d6c3c3f081f5,64'hdfffffff20000001,
64'h585bda2e086ebc26,64'h0000003fffbfffc0,64'h80b6b6221f840fa4,64'h0000000000000001
};
  //------------------------
  // 64
  //------------------------
  localparam [2*64-1:0][63:0] NTT_GF64_BWD_N64_PHI_L = {
64'h000001fffdfffe00,64'h0000000000000008,64'h00000fffeffff000,64'h0000000000000040,
64'h00007fff7fff8000,64'h0000000000000200,64'h0003fffbfffc0000,64'h0000000000001000,
64'h001fffdfffe00000,64'h0000000000008000,64'h00fffeffff000000,64'h0000000000040000,
64'h07fff7fff8000000,64'h0000000000200000,64'h3fffbfffc0000000,64'h0000000001000000,
64'hfffdfffeffffffff,64'h0000000008000000,64'hffeffffefffffff1,64'h0000000040000000,
64'hff7ffffeffffff81,64'h0000000200000000,64'hfbfffffefffffc01,64'h0000001000000000,
64'hdffffffeffffe001,64'h0000008000000000,64'hfffffffdffff0002,64'h0000040000000000,
64'hfffffff6fff80009,64'h0000200000000000,64'hffffffbeffc00041,64'h0001000000000000,
64'hfffffdfefe000201,64'h0008000000000000,64'hffffeffef0001001,64'h0040000000000000,
64'hffff7ffe80008001,64'h0200000000000000,64'hfffbfffb00040001,64'h1000000000000000,
64'hffdfffdf00200001,64'h8000000000000000,64'hfefffeff01000001,64'h00000003fffffffc,
64'hf7fff7ff08000001,64'h0000001fffffffe0,64'hbfffbfff40000001,64'h000000ffffffff00,
64'hfffdffff00000003,64'h000007fffffff800,64'hffefffff00000011,64'h00003fffffffc000,
64'hff7fffff00000081,64'h0001fffffffe0000,64'hfbffffff00000401,64'h000ffffffff00000,
64'hdfffffff00002001,64'h007fffffff800000,64'hfffffffe00010002,64'h03fffffffc000000,
64'hfffffff700080009,64'h1fffffffe0000000,64'hffffffbf00400041,64'hffffffff00000000,
64'hfffffdff02000201,64'hfffffffefffffff9,64'hffffefff10001001,64'hfffffffeffffffc1,
64'hffff7fff80008001,64'hfffffffefffffe01,64'hfffc000300040001,64'hfffffffefffff001,
64'hffe0001f00200001,64'hfffffffeffff8001,64'hff0000ff01000001,64'hfffffffefffc0001,
64'hf80007ff08000001,64'hfffffffeffe00001,64'hc0003fff40000001,64'hfffffffeff000001,
64'h0002000000000002,64'hfffffffef8000001,64'h0010000000000010,64'hfffffffec0000001,
64'h0080000000000080,64'hfffffffd00000001,64'h0400000000000400,64'hffffffef00000001,
64'h2000000000002000,64'hffffff7f00000001,64'h000000010000ffff,64'hfffffbff00000001,
64'h000000080007fff8,64'hffffdfff00000001,64'h00000040003fffc0,64'hfffeffff00000001,
64'h0000020001fffe00,64'hfff7ffff00000001,64'h000010000ffff000,64'hffbfffff00000001,
64'h000080007fff8000,64'hfdffffff00000001,64'h00040003fffc0000,64'hefffffff00000001,
64'h0020001fffe00000,64'h7fffffff00000001,64'h010000ffff000000,64'hfffffffb00000005,
64'h080007fff8000000,64'hffffffdf00000021,64'h40003fffc0000000,64'hfffffeff00000101,
64'h0001fffffffffffe,64'hfffff7ff00000801,64'h000ffffffffffff0,64'hffffbfff00004001,
64'h007fffffffffff80,64'hfffdffff00020001,64'h03fffffffffffc00,64'hffefffff00100001,
64'h1fffffffffffe000,64'hff7fffff00800001,64'h00000000fffeffff,64'hfbffffff04000001,
64'h00000007fff7fff8,64'hdfffffff20000001,64'h0000003fffbfffc0,64'h0000000000000001
};
  //------------------------
  // 32
  //------------------------
  localparam [2*32-1:0][63:0] NTT_GF64_BWD_N32_PHI_L = {
64'h0000000000000008,64'h0000000000000040,64'h0000000000000200,64'h0000000000001000,
64'h0000000000008000,64'h0000000000040000,64'h0000000000200000,64'h0000000001000000,
64'h0000000008000000,64'h0000000040000000,64'h0000000200000000,64'h0000001000000000,
64'h0000008000000000,64'h0000040000000000,64'h0000200000000000,64'h0001000000000000,
64'h0008000000000000,64'h0040000000000000,64'h0200000000000000,64'h1000000000000000,
64'h8000000000000000,64'h00000003fffffffc,64'h0000001fffffffe0,64'h000000ffffffff00,
64'h000007fffffff800,64'h00003fffffffc000,64'h0001fffffffe0000,64'h000ffffffff00000,
64'h007fffffff800000,64'h03fffffffc000000,64'h1fffffffe0000000,64'hffffffff00000000,
64'hfffffffefffffff9,64'hfffffffeffffffc1,64'hfffffffefffffe01,64'hfffffffefffff001,
64'hfffffffeffff8001,64'hfffffffefffc0001,64'hfffffffeffe00001,64'hfffffffeff000001,
64'hfffffffef8000001,64'hfffffffec0000001,64'hfffffffd00000001,64'hffffffef00000001,
64'hffffff7f00000001,64'hfffffbff00000001,64'hffffdfff00000001,64'hfffeffff00000001,
64'hfff7ffff00000001,64'hffbfffff00000001,64'hfdffffff00000001,64'hefffffff00000001,
64'h7fffffff00000001,64'hfffffffb00000005,64'hffffffdf00000021,64'hfffffeff00000101,
64'hfffff7ff00000801,64'hffffbfff00004001,64'hfffdffff00020001,64'hffefffff00100001,
64'hff7fffff00800001,64'hfbffffff04000001,64'hdfffffff20000001,64'h0000000000000001
};
  //------------------------
  // 16
  //------------------------
  localparam [2*16-1:0][63:0] NTT_GF64_BWD_N16_PHI_L = {
64'h0000000000000040,64'h0000000000001000,64'h0000000000040000,64'h0000000001000000,
64'h0000000040000000,64'h0000001000000000,64'h0000040000000000,64'h0001000000000000,
64'h0040000000000000,64'h1000000000000000,64'h00000003fffffffc,64'h000000ffffffff00,
64'h00003fffffffc000,64'h000ffffffff00000,64'h03fffffffc000000,64'hffffffff00000000,
64'hfffffffeffffffc1,64'hfffffffefffff001,64'hfffffffefffc0001,64'hfffffffeff000001,
64'hfffffffec0000001,64'hffffffef00000001,64'hfffffbff00000001,64'hfffeffff00000001,
64'hffbfffff00000001,64'hefffffff00000001,64'hfffffffb00000005,64'hfffffeff00000101,
64'hffffbfff00004001,64'hffefffff00100001,64'hfbffffff04000001,64'h0000000000000001
};
  //------------------------
  // 8
  //------------------------
  localparam [2*8-1:0][63:0] NTT_GF64_BWD_N8_PHI_L = {
64'h0000000000001000,64'h0000000001000000,64'h0000001000000000,64'h0001000000000000,
64'h1000000000000000,64'h000000ffffffff00,64'h000ffffffff00000,64'hffffffff00000000,
64'hfffffffefffff001,64'hfffffffeff000001,64'hffffffef00000001,64'hfffeffff00000001,
64'hefffffff00000001,64'hfffffeff00000101,64'hffefffff00100001,64'h0000000000000001
};
  //------------------------
  // 4
  //------------------------
  localparam [2*4-1:0][63:0] NTT_GF64_BWD_N4_PHI_L = {
64'h0000000001000000,64'h0001000000000000,64'h000000ffffffff00,64'hffffffff00000000,
64'hfffffffeff000001,64'hfffeffff00000001,64'hfffffeff00000101,64'h0000000000000001
};

  //========================
  // NTT backward with div 1/N
  //========================
  //------------------------
  // 2048
  //------------------------
  localparam [2*2048-1:0][63:0] NTT_GF64_BWD_WDIV_N2048_PHI_L = {
64'h197309d889c9a00b,64'h030f4b22afbccf85,64'h7a5c0850fca5dae7,64'ha8c7b40b550e189f,
64'h39a8014de318bf1a,64'hf84069b87c7158a1,64'h9a6f702a47793880,64'h55f9087dd6728c17,
64'h2653648b9aca776b,64'h96bfeb83763604e6,64'h8b0355af4298a8e1,64'h214735f58c465163,
64'ha88614e450d3cae7,64'hbecadd83091f60a1,64'h30804f6245d269bc,64'hda585bd954086ebd,
64'hda815a870160d25a,64'hdaae61c6df8f42f0,64'h0094a678f8ec1661,64'h6b817fb2f1af13a5,
64'hcea9a8b27ab0509e,64'h848743e4022bde2c,64'h0776f3d907a932c4,64'h7a4b539d96a7c922,
64'hb6cceb510e610f9c,64'hed0e4676e0541588,64'h12ee4830e85a03de,64'hd4897a64274f5176,
64'h29a8b8e589433675,64'hc4e614a1c6e8d04d,64'h3cedaf0525e1493c,64'h3fffffffffffc000,
64'he1f99c7870df1f01,64'h343971c45dd0cf37,64'ha8c7c9442f2e4818,64'h0435911517b83abe,
64'h9544b20b4af2803d,64'h6fc7dc8a5c6bcddb,64'h9cad2d792fe38a52,64'he8bf5629fb82c865,
64'h7d6c99faee94b994,64'h63efdef1494caceb,64'hd1b688ec0718e627,64'ha147aaae1f33dd54,
64'hdda318ee7f917589,64'h37316c05eb014da9,64'hdfe6d22be2eec414,64'h5c80b6b5c61f8410,
64'hb1ecedf0895b40b3,64'h8f116300a66bef05,64'he639c0843c87755c,64'hf76ce80155b0531d,
64'hfa0e866f11aab25d,64'h8eaef0b242c4ee84,64'ha04747a337c1b3d9,64'h13705cd1d6bb177a,
64'h1e94da9c6d77bfba,64'hb890496d2d221ecd,64'h52112b41b38dbec0,64'hd4ab38be64115ea7,
64'hbb0711cd3e749c60,64'h8c88faabc9bfee9c,64'hb7ccd994ea895913,64'hfeffffff01000001,
64'hcb984ec44e4d0058,64'h187a59157de67c28,64'hd2e0428ae52ed735,64'h463da05fa870c4f3,
64'hcd400a7018c5f8cf,64'hc2034dcae38ac501,64'hd37b81563bc9c3fc,64'hafc843f0b39460b6,
64'h329b245dd653bb57,64'hb5ff5c1fb1b0272c,64'h581aad7e14c54704,64'h0a39afad62328b17,
64'h4430a727869e5733,64'hf656ec1d48fb0503,64'h84027b132e934ddf,64'hd2c2ded0a04375e2,
64'hd40ad43e0b0692ca,64'hd5730e3cfc7a177a,64'h04a533c7c760b308,64'h5c0bfd9a8d789d25,
64'h754d4599d58284ea,64'h243a1f24115ef15c,64'h3bb79ec83d499620,64'hd25a9cefb53e490d,
64'hb6675a8d73087cdb,64'h687233be02a0ac39,64'h9772418742d01ef0,64'ha44bd3273a7a8baa,
64'h4d45c72d4a19b3a7,64'h2730a51437468262,64'he76d782a2f0a49df,64'h00000001fffdfffe,
64'h0fcce3ca86f8f801,64'ha1cb8e23ee8679b7,64'h463e4a26797240bb,64'h21ac88a8bdc1d5f0,
64'haa25905e579401e4,64'h7e3ee455e35e6ed5,64'he5696bcd7f1c528c,64'h45fab156dc164321,
64'heb64cfda74a5cc9d,64'h1f7ef78d4a656755,64'h8db4476638c73132,64'h0a3d5575f99eea9b,
64'hed18c779fc8bac42,64'hb98b6030580a6d47,64'hff3691651776209a,64'he405b5b030fc207e,
64'h8f676f894ada0593,64'h788b1809335f7824,64'h31ce0428e43baad9,64'hbb674011ad8298e1,
64'hd074337f8d5592e1,64'h757785961627741c,64'h023a3d1ebe0d9ec3,64'h9b82e68eb5d8bbd0,
64'hf4a6d4e36bbdfdd0,64'hc4824b6e6910f663,64'h90895a0f9c6df5fe,64'ha559c5f9208af532,
64'hd8388e6ef3a4e2fb,64'h6447d5624dff74dc,64'hbe66ccac544ac893,64'hf7ffffff08000001,
64'h5cc27628726802ba,64'hc3d2c8abef33e140,64'h9702145d2976b9a2,64'h31ed02ff43862796,
64'h6a005386c62fc672,64'h101a6e5d1c562802,64'h9bdc0ab7de4e1fda,64'h7e421f8a9ca305ab,
64'h94d922efb29ddab7,64'haffae1028d81395b,64'hc0d56bf2a62a381e,64'h51cd7d6b119458b8,
64'h2185393e34f2b996,64'hb2b760f147d82811,64'h2013d89d749a6ef4,64'h9616f68b021baf0a,
64'ha056a1f65834964a,64'hab9871ede3d0bbca,64'h25299e3e3b059840,64'he05fecd66bc4e926,
64'haa6a2cd1ac14274d,64'h21d0f9218af78adf,64'hddbcf642ea4cb0ff,64'h92d4e783a9f24862,
64'hb33ad4709843e6d3,64'h43919df3150561c5,64'hbb920c3e1680f77c,64'h225e993ed3d45d4b,
64'h6a2e396c50cd9d36,64'h398528a2ba34130f,64'h3b6bc15878524ef1,64'h0000000fffeffff0,
64'h7e671e5437c7c008,64'h0e5c71247433cdb3,64'h31f25135cb9205d6,64'h0d644546ee0eaf7f,
64'h512c82f7bca00f1b,64'hf1f722b21af376a5,64'h2b4b5e72f8e29459,64'h2fd58ab8e0b21906,
64'h5b267edaa52e64e1,64'hfbf7bc6a532b3aa8,64'h6da23b35c639898c,64'h51eaabafccf754d8,
64'h68c63bd6e45d6209,64'hcc5b0187c0536a33,64'hf9b48b2fbbb104c9,64'h202dad8887e103e9,
64'h7b3b7c4e56d02c94,64'hc458c04c9afbc11d,64'h8e70214821dd56c7,64'hdb3a00926c14c703,
64'h83a19c026aac9702,64'habbc2cb3b13ba0dd,64'h11d1e8f5f06cf618,64'hdc173479aec5de7c,
64'ha536a7225defee79,64'h24125b794887b312,64'h844ad080e36fafec,64'h2ace2fce0457a98b,
64'hc1c4737d9d2717d2,64'h223eab156ffba6dd,64'hf3366567a2564493,64'hbfffffff40000001,
64'he613b145934015ce,64'h1e964565799f09fa,64'hb810a2ed4bb5cd0c,64'h8f6817fb1c313caf,
64'h50029c39317e338d,64'h80d372e8e2b14010,64'hdee055c2f270fecc,64'hf210fc57e5182d55,
64'ha6c9178194eed5b4,64'h7fd708196c09cad3,64'h06ab5f9b3151c0ea,64'h8e6beb5a8ca2c5be,
64'h0c29c9f2a795ccaf,64'h95bb078f3ec14083,64'h009ec4eca4d3779f,64'hb0b7b45c10dd784c,
64'h02b50fb7c1a4b24b,64'h5cc38f741e85de4b,64'h294cf1f2d82cc1ff,64'h02ff66ba5e274929,
64'h5351669260a13a63,64'h0e87c90d57bc56f7,64'hede7b21d526587f2,64'h96a73c214f92430c,
64'h99d6a389c21f3693,64'h1c8cef9aa82b0e26,64'hdc9061f5b407bbdb,64'h12f4c9f79ea2ea57,
64'h5171cb65866ce9ad,64'hcc294516d1a09877,64'hdb5e0ac4c2927787,64'h0000007fff7fff80,
64'hf338f2a4be3e003d,64'h72e38923a19e6d98,64'h8f9289af5c902eaf,64'h6b222a3770757bf8,
64'h896417bfe50078d6,64'h8fb91597d79bb521,64'h5a5af398c714a2c7,64'h7eac55c80590c82f,
64'hd933f6d729732706,64'hdfbde3599959d539,64'h6d11d9b131cc4c5d,64'h8f555d8067baa6be,
64'h4631deba22eb1045,64'h62d80c44029b5192,64'hcda45984dd882641,64'h016d6c453f081f47,
64'hd9dbe275b681649d,64'h22c6026ad7de08e2,64'h73810a450eeab634,64'hd9d0049960a63812,
64'h1d0ce0175564b80c,64'h5de165a289dd06e3,64'h8e8f47af8367b0c0,64'he0b9a3d3762ef3da,
64'h29b53917ef7f73c3,64'h2092dbcb443d988f,64'h2256840b1b7d7f5c,64'h56717e7122bd4c57,
64'h0e239bf2e938be8a,64'h11f558ac7fdd36e7,64'h99b32b4412b22491,64'h0000000000000002,
64'h309d8a339a00ae69,64'hf4b22b2bccf84fd0,64'hc085176f5dae685b,64'h7b40bfdce189e574,
64'h8014e1cb8bf19c66,64'h069b974b158a007c,64'hf702ae1d9387f65a,64'h9087e2c628c16aa1,
64'h3648bc11a776ad9b,64'hfeb840ce604e5695,64'h355afcd98a8e0750,64'h735f5ad865162dec,
64'h614e4f953cae6578,64'hadd83c7df60a0414,64'h04f62765269bbcf8,64'h85bda2e586ebc25b,
64'h15a87dbe0d259258,64'he61c7ba2f42ef256,64'h4a678f97c1660ff7,64'h17fb35d2f13a4948,
64'h9a8b34950509d316,64'h743e486abde2b7b8,64'h6f3d90f1932c3f89,64'hb539e10e7c92185c,
64'hceb51c5210f9b494,64'he4677cd541587130,64'he4830fb3a03dded2,64'h97a64fbcf51752b8,
64'h8b8e5b2e33674d66,64'h614a28bc8d04c3b2,64'hdaf0562c1493bc32,64'h000003fffbfffc00,
64'h99c7952cf1f001e1,64'h971c49200cf36cbd,64'h7c944d7ee4817574,64'h591151be83abdfbd,
64'h4b20be032803c6ac,64'h7dc8acc2bcdda904,64'hd2d79cc838a51636,64'hf562ae432c864175,
64'hc99fb6bf4b99382a,64'hfdef1ad2cacea9c2,64'h688ecd8c8e6262e5,64'h7aaaec073dd535ec,
64'h318ef5d317588226,64'h16c0622314da8c8d,64'h6d22cc2cec413202,64'h0b6b6229f840fa38,
64'hcedf13b3b40b24e2,64'h16301357bef0470f,64'h9c08522b7755b19d,64'hce8024d10531c08a,
64'he86700baab25c060,64'hef0b2d164ee83716,64'h747a3d801b3d85fc,64'h05cd1ea2b1779ec9,
64'h4da9c8c07bfb9e17,64'h0496de5b21ecc477,64'h12b42059dbebfadf,64'hb38bf38b15ea62b6,
64'h711cdf9749c5f450,64'h8faac563fee9b738,64'hcd995a2495912484,64'h0000000000000010,
64'h84ec519dd0057347,64'ha591596567c27e79,64'h0428bb80ed7342d2,64'hda05feea0c4f2b9d,
64'h00a70e605f8ce32c,64'h34dcba58ac5003e0,64'hb81570f39c3fb2c9,64'h843f1635460b5504,
64'hb245e08e3bb56cd7,64'hf5c2067a0272b4a1,64'haad7e6cd54703a7f,64'h9afad6c628b16f5d,
64'h0a727cace5732bbd,64'h6ec1e3f4b050209b,64'h27b13b2934dde7c0,64'h2ded1730375e12d4,
64'had43edf0692c92c0,64'h30e3dd1ea17792a9,64'h533c7cc00b307fb6,64'hbfd9ae9789d24a40,
64'hd459a4ac284e98ac,64'ha1f24358ef15bdbd,64'h79ec878f9961fc45,64'ha9cf0878e490c2db,
64'h75a8e29687cda49a,64'h233be6b10ac38979,64'h24187da401eef689,64'hbd327deba8ba95bc,
64'h5c72d9759b3a6b2c,64'h0a5145e768261d8d,64'hd782b166a49de18a,64'h00001fffdfffe000,
64'hce3ca96b8f800f04,64'hb8e24904679b65e4,64'he4a26bfa240bab9d,64'hc88a8df61d5efde6,
64'h5905f01b401e355e,64'hee456618e6ed481d,64'h96bce647c528b1aa,64'hab15722064320ba1,
64'h4cfdb6005cc9c14a,64'hef78d69d56754e09,64'h44766c6773131725,64'hd557603ceea9af5d,
64'h8c77ae99bac4112f,64'hb6031118a6d46468,64'h6916616a6209900d,64'h5b5b114fc207d1c0,
64'h76f89da3a059270a,64'hb1809abdf7823878,64'he042915fbaad8ce4,64'h7401268e298e044a,
64'h433805dc592e02f9,64'h785968b97741b8a9,64'ha3d1ec03d9ec2fdd,64'h2e68f5158bbcf648,
64'h6d4e4605dfdcf0b6,64'h24b6f2d90f6623b8,64'h95a102cedf5fd6f8,64'h9c5f9c5daf5315ab,
64'h88e6fcbd4e2fa27d,64'h7d562b23f74db9bc,64'h6ccad12aac89241a,64'h0000000000000080,
64'h27628cf2802b9a34,64'h2c8acb303e13f3c3,64'h2145dc076b9a1690,64'hd02ff75662795ce2,
64'h05387302fc671960,64'ha6e5d2c662801eff,64'hc0ab87a1e1fd9643,64'h21f8b1ae305aa81c,
64'h922f0476ddab66b3,64'hae1033d71395a501,64'h56bf366fa381d3f3,64'hd7d6b635458b7ae4,
64'h5393e5672b995de8,64'h760f1fa8828104d5,64'h3d89d94aa6ef3dff,64'h6f68b982baf0969f,
64'h6a1f6f88496495fb,64'h871ee8f60bbc9547,64'h99e3e6025983fdae,64'hfecd74c14e9251fb,
64'ha2cd25674274c55a,64'h0f921acc78adede3,64'hcf643c7fcb0fe225,64'h4e7843cc248616d3,
64'had4714b73e6d24cd,64'h19df3589561c4bc7,64'h20c3ed210f77b447,64'he993ef6245d4addb,
64'he396cbaed9d3595e,64'h528a2f3b4130ec68,64'hbc158b3b24ef0c4a,64'h0000fffeffff0000,
64'h71e54b627c00781a,64'hc71248283cdb2f1b,64'h25135fd8205d5ce1,64'h44546fb6eaf7ef2a,
64'hc82f80dc00f1aaee,64'h722b30ce376a40e1,64'hb5e7324229458d4c,64'h58ab910821905d03,
64'h67edb004e64e0a4e,64'h7bc6b4f1b3aa7041,64'h23b3633d9898b926,64'haabb01ed754d7ae2,
64'h63bd74d1d6208974,64'hb01888ca36a3233b,64'h48b30b56104c8065,64'hdad88a80103e8dfe,
64'hb7c4ed2002c9384d,64'h8c04d5f4bc11c3bb,64'h02148b04d56c6719,64'ha00934744c70224d,
64'h19c02ee4c97017c6,64'hc2cb45ceba0dc545,64'h1e8f6023cf617ee3,64'h7347a8ad5de7b23f,
64'h6a723031fee785ad,64'h25b796c97b311dbf,64'had08167afafeb7bc,64'he2fce2f17a98ad54,
64'h4737e5ee717d13e4,64'heab15922ba6dcddd,64'h66568958644920cd,64'h0000000000000400,
64'h3b146795015cd19f,64'h64565982f09f9e17,64'h0a2ee03c5cd0b47f,64'h817fbab913cae70a,
64'h29c39817e338cb00,64'h372e96381400f7f3,64'h055c3d150fecb212,64'h0fc58d7282d540df,
64'h917823baed5b3594,64'h70819ebd9cad2803,64'hb5f9b37f1c0e9f96,64'hbeb5b1b02c5bd71a,
64'h9c9f2b3b5ccaef3e,64'hb078fd47140826a5,64'hec4eca563779eff7,64'h7b45cc18d784b4f5,
64'h50fb7c454b24afd5,64'h38f747b45de4aa34,64'hcf1f3016cc1fed6c,64'hf66ba61174928fd1,
64'h16692b3f13a62acb,64'h7c90d663c56f6f18,64'h7b21e404587f1122,64'h73c21e632430b696,
64'h6a38a5bef3692663,64'hcef9ac4ab0e25e38,64'h061f69097bbda237,64'h4c9f7b192ea56ed1,
64'h1cb65d7dce9acae9,64'h945179dc0987633e,64'he0ac59de2778624b,64'h0007fff7fff80000,
64'h8f2a5b16e003c0cd,64'h38924147e6d978d2,64'h289afec202eae707,64'h22a37db957bf794e,
64'h417c06e6078d576a,64'h91598674bb520705,64'haf3992164a2c6a5b,64'hc55c88430c82e816,
64'h3f6d802a3270526d,64'hde35a7909d538205,64'h1d9b19edc4c5c92f,64'h55d80f70aa6bd70b,
64'h1deba691b1044b9d,64'h80c44656b51919d3,64'h45985ab282640326,64'hd6c4540681f46fea,
64'hbe2769051649c263,64'h6026afa9e08e1dd4,64'h10a45826ab6338c8,64'h0049a3a763811263,
64'hce0177264b80be30,64'h165a2e7bd06e2a22,64'hf47b011e7b0bf718,64'h9a3d456def3d91f5,
64'h53918192f73c2d65,64'h2dbcb64cd988edf7,64'h6840b3dcd7f5bddb,64'h17e71792d4c56a99,
64'h39bf2f758be89f1e,64'h558ac91cd36e6ee1,64'h32b44ac622490665,64'h0000000000002000,
64'hd8a33ca90ae68cf7,64'h22b2cc1a84fcf0b5,64'h517701e2e685a3f8,64'h0bfdd5cc9e57384c,
64'h4e1cc0c019c657ff,64'hb974b1c1a007bf97,64'h2ae1e8a87f659090,64'h7e2c6b9416aa06f8,
64'h8bc11ddb6ad9ac9c,64'h840cf5efe5694015,64'hafcd9bfde074fcab,64'hf5ad8d8662deb8cb,
64'he4f959dee65779ec,64'h83c7ea3da0413523,64'h627652b8bbcf7fb1,64'hda2e60c9bc25a7a5,
64'h87dbe22c59257ea6,64'hc7ba3da3ef25519f,64'h78f980bc60ff6b5a,64'hb35d3092a4947e81,
64'hb34959f89d315658,64'he486b3212b7b78bd,64'hd90f2025c3f8890d,64'h9e10f31c2185b4ad,
64'h51c52dfa9b493315,64'h77cd625b8712f1ba,64'h30fb484bdded11b8,64'h64fbd8cb752b7686,
64'he5b2ebee74d65748,64'ha28bcee44c3b19ec,64'h0562cef83bc31251,64'h003fffbfffc00000,
64'h7952d8bb001e0664,64'hc4920a4036cbc68f,64'h44d7f61117573837,64'h151bedcbbdfbca6f,
64'h0be037323c6abb4e,64'h8acc33a9da903824,64'h79cc90b7516352d3,64'h2ae4421e641740aa,
64'hfb6c015293829367,64'hf1ad3c8aea9c1022,64'hecd8cf6e262e4978,64'haec07b87535eb856,
64'hef5d348d88225ce8,64'h062232b9a8c8ce94,64'h2cc2d5961320192e,64'hb622a03a0fa37f4a,
64'hf13b482db24e1313,64'h01357d520470ee9d,64'h8522c1355b19c640,64'h024d1d3b1c089318,
64'h700bb9385c05f17a,64'hb2d173de83715110,64'ha3d808fad85fb8b9,64'hd1ea2b7379ec8fa4,
64'h9c8c0c99b9e16b26,64'h6de5b267cc476fb7,64'h42059ee9bfadeed5,64'hbf38bc96a62b54c8,
64'hcdf97bad5f44f8ef,64'hac5648e89b737706,64'h95a2563212483327,64'h0000000000010000,
64'hc519e54e573467b2,64'h159660d527e785a7,64'h8bb80f19342d1fbe,64'h5feeae64f2b9c260,
64'h70e60602ce32bff6,64'hcba58e12003dfcb3,64'h570f4544fb2c847f,64'hf1635ca3b55037bd,
64'h5e08eedf56cd64dc,64'h2067af832b4a00a4,64'h7e6cdff403a7e553,64'had6c6c3a16f5c651,
64'h27cacefe32bbcf59,64'h1e3f51f10209a914,64'h13b295c8de7bfd85,64'hd1730653e12d3d22,
64'h3edf1166c92bf52c,64'h3dd1ed25792a8cf2,64'hc7cc05e607fb5acd,64'h9ae9849a24a3f403,
64'h9a4acfc9e98ab2bb,64'h243599105bdbc5e1,64'hc87901341fc44862,64'hf08798e50c2da564,
64'h8e296fd6da4998a6,64'hbe6b12df38978dcd,64'h87da425fef688dbf,64'h27dec65ea95bb42d,
64'h2d975f7aa6b2ba39,64'h145e772761d8cf5b,64'h2b1677c1de189288,64'h01fffdfffe000000,
64'hca96c5db00f0331d,64'h24905207b65e3472,64'h26bfb08abab9c1b6,64'ha8df6e5defde5378,
64'h5f01b991e355da70,64'h56619d52d481c11c,64'hce6485bd8b1a9695,64'h572210f420ba054f,
64'hdb600a9b9c149b31,64'h8d69e45e54e08109,64'h66c67b7831724bb9,64'h7603dc3f9af5c2ab,
64'h7ae9a4734112e739,64'h311195cd464674a0,64'h6616acb19900c96f,64'hb11501d57d1bfa4b,
64'h89da417492709891,64'h09abea90238774e8,64'h291609aed8ce31fc,64'h1268e9d8e04498c0,
64'h805dc9c5e02f8bcd,64'h968b9ef91b8a887b,64'h1ec047dbc2fdc5c3,64'h8f515ba1cf647d1a,
64'he46064d1cf0b592c,64'h6f2d9341623b7db5,64'h102cf74ffd6f76a6,64'hf9c5e4ba315aa63b,
64'h6fcbdd70fa27c772,64'h62b24749db9bb82b,64'had12b19492419934,64'h0000000000080000,
64'h28cf2a78b9a33d8a,64'hacb306a93f3c2d38,64'h5dc078cda168fdec,64'hff75732995ce12fe,
64'h873030197195ffad,64'h5d2c709601efe592,64'hb87a2a29d96423f6,64'h8b1ae524aa81bde1,
64'hf04776fcb66b26de,64'h033d7c1a5a50051f,64'hf366ffa31d3f2a95,64'h6b6361d5b7ae3283,
64'h3e5677f295de7ac7,64'hf1fa8f88104d48a0,64'h9d94ae46f3dfec28,64'h8b9832a50969e90a,
64'hf6f88b37495fa95f,64'hee8f692cc954678f,64'h3e602f363fdad662,64'hd74c24d5251fa014,
64'hd2567e534c5595d4,64'h21acc883dede2f07,64'h43c809a6fe22430a,64'h843cc72f616d2b19,
64'h714b7ebad24cc52c,64'hf35896fec4bc6e63,64'h3ed213037b446df4,64'h3ef632f64adda167,
64'h6cbafbd63595d1c7,64'ha2f3b93b0ec67ad8,64'h58b3be0ff0c4943f,64'h0fffeffff0000000,
64'h54b62ede078198e2,64'h2482903eb2f1a38f,64'h35fd8456d5ce0daf,64'h46fb72f47ef29bbb,
64'hf80dcc911aaed37e,64'hb30cea98a40e08de,64'h73242df258d4b4a2,64'hb91087a305d02a76,
64'hdb0054e2e0a4d982,64'h6b4f22f6a7040844,64'h3633dbc48b925dc5,64'hb01ee1ffd7ae1555,
64'hd74d239d089739c5,64'h888cae6b3233a4ff,64'h30b5658fc8064b75,64'h88a80eb0e8dfd253,
64'h4ed20ba89384c484,64'h4d5f54811c3ba740,64'h48b04d77c6718fdf,64'h93474ec70224c600,
64'h02ee4e33017c5e64,64'hb45cf7ccdc5443d4,64'hf6023ede17ee2e18,64'h7a8add127b23e8cc,
64'h23032695785ac959,64'h796c9a0e11dbeda5,64'h8167ba7feb7bb530,64'hce2f25d88ad531d1,
64'h7e5eeb8ad13e3b8d,64'h15923a51dcddc155,64'h68958ca9920cc99b,64'h0000000000400000,
64'h467953c6cd19ec4f,64'h6598354ef9e169bb,64'hee03c66f0b47ef5e,64'hfbab9953ae7097e9,
64'h398180cf8caffd64,64'he96384b20f7f2c8e,64'hc3d15153cb211fab,64'h58d72929540def04,
64'h823bb7ecb35936e9,64'h19ebe0d2d28028f8,64'h9b37fd1fe9f954a1,64'h5b1b0eb0bd719415,
64'hf2b3bf95aef3d637,64'h8fd47c47826a44f9,64'heca5723b9eff613c,64'h5cc1952c4b4f484c,
64'hb7c459c14afd4af1,64'h747b496d4aa33c71,64'hf30179b2fed6b30f,64'hba6126af28fd009a,
64'h92b3f2a062acae9a,64'h0d66441ff6f17837,64'h1e404d39f112184e,64'h21e6397f0b6958c4,
64'h8a5bf5d99266295d,64'h9ac4b7fd25e37311,64'hf690981cda236f9f,64'hf7b197b356ed0b37,
64'h65d7deb4acae8e35,64'h179dc9dd7633d6bb,64'hc59df0818624a1f6,64'h7fff7fff80000000,
64'ha5b176f23c0cc70e,64'h241481f6978d1c77,64'hafec22b7ae706d77,64'h37db97a5f794ddd6,
64'hc06e648fd5769be9,64'h986754ca207046eb,64'h99216f95c6a5a50d,64'hc8843d1d2e8153ab,
64'hd802a71d0526cc0a,64'h5a7917b83820421d,64'hb19ede255c92ee27,64'h80f71003bd70aaa3,
64'hba691cee44b9ce22,64'h4465735d919d27f4,64'h85ab2c7f40325ba7,64'h4540758b46fe9294,
64'h76905d469c26241e,64'h6afaa40ae1dd39fe,64'h45826bc0338c7ef6,64'h9a3a763c11262ffc,
64'h177271980be2f320,64'ha2e7be6be2a21e9b,64'hb011f6f7bf7170b9,64'hd456e896d91f465d,
64'h181934acc2d64ac7,64'hcb64d0738edf6d25,64'h0b3dd4035bdda97c,64'h71792eca56a98e82,
64'hf2f75c5989f1dc65,64'hac91d28ee6ee0aa8,64'h44ac654f90664cd5,64'h0000000002000000,
64'h33ca9e3868cf6276,64'h2cc1aa7acf0b4dd5,64'h701e337f5a3f7ae9,64'hdd5ccaa47384bf41,
64'hcc0c067d657feb1f,64'h4b1c25977bf96469,64'h1e8a8aa45908fd52,64'hc6b9494ca06f781e,
64'h11ddbf699ac9b744,64'hcf5f0696940147c0,64'hd9bfe9034fcaa504,64'hd8d87587eb8ca0a6,
64'h959dfcb4779eb1b1,64'h7ea3e240135227c4,64'h652b91e3f7fb09d9,64'he60ca9645a7a425e,
64'hbe22ce0f57ea5783,64'ha3da4b6d5519e385,64'h980bcd9ef6b59871,64'hd309357e47e804cb,
64'h959f9507156574cc,64'h6b3220ffb78bc1b8,64'hf20269cf8890c270,64'h0f31cbf95b4ac61f,
64'h52dfaed093314ae4,64'hd625bfed2f1b9884,64'hb484c0edd11b7cf1,64'hbd8cbda1b76859b1,
64'h2ebef5a8657471a5,64'hbcee4eebb19eb5d8,64'h2cef841231250faa,64'hfffbfffefffffffd,
64'h2d8bb796e066386b,64'h20a40fb5bc68e3b7,64'h7f6115c273836bb3,64'hbedcbd30bca6eeaf,
64'h03732484abb4df42,64'hc33aa65503823754,64'hc90b7cb2352d2864,64'h4421e8ef740a9d52,
64'hc01538ee2936604a,64'hd3c8bdc3c10210e6,64'h8cf6f12fe4977133,64'h07b88021eb855514,
64'hd348e77725ce710b,64'h232b9aee8ce93f9e,64'h2d5963fe0192dd34,64'h2a03ac5c37f4949e,
64'hb482ea37e13120ed,64'h57d5205a0ee9cfed,64'h2c135e039c63f7ae,64'hd1d3b1e489317fdc,
64'hbb938cc05f179900,64'h173df3641510f4d3,64'h808fb7c2fb8b85c3,64'ha2b744bcc8fa32e2,
64'hc0c9a56616b25638,64'h5b2683a276fb6922,64'h59eea01adeed4be0,64'h8bc97655b54c740d,
64'h97bae2d34f8ee321,64'h648e947c3770553b,64'h25632a7e833266a6,64'h0000000010000000,
64'h9e54f1c4467b13af,64'h660d53d7785a6ea7,64'h80f19bfdd1fbd745,64'heae655299c25fa02,
64'h606033f12bff58f2,64'h58e12cbddfcb2346,64'hf4545522c847ea90,64'h35ca4a6b037bc0ea,
64'h8eedfb4cd64dba20,64'h7af834baa00a3dfa,64'hcdff48207e55281a,64'hc6c3ac455c65052a,
64'hacefe5a7bcf58d84,64'hf51f12039a913e1d,64'h295c8f22bfd84ec5,64'h30654b29d3d212e9,
64'hf116707fbf52bc13,64'h1ed25b6fa8cf1c23,64'hc05e6cfbb5acc384,64'h9849abf83f402652,
64'hacfca83cab2ba65c,64'h59910800bc5e0dbd,64'h90134e8344861379,64'h798e5fcada5630f8,
64'h96fd7686998a571e,64'hb12dff6f78dcc41a,64'ha426077388dbe783,64'hec65ed12bb42cd83,
64'h75f7ad442ba38d27,64'he77277628cf5aebb,64'h677c209289287d4f,64'hffdffffeffffffe1,
64'h6c5dbcb80331c357,64'h05207daee3471db7,64'hfb08ae169c1b5d95,64'hf6e5e98ae5377573,
64'h1b9924255da6fa10,64'h19d532ae1c11ba9a,64'h485be597a969431a,64'h210f477da054ea8e,
64'h00a9c77749b3024a,64'h9e45ee240810872a,64'h67b7898324bb8994,64'h3dc4010f5c2aa8a0,
64'h9a473bbf2e738852,64'h195cd7756749fcef,64'h6acb1ff10c96e99f,64'h501d62e2bfa4a4ef,
64'ha41751c409890763,64'hbea902d2774e7f66,64'h609af01de31fbd6f,64'h8e9d8f2a498bfeda,
64'hdc9c6607f8bcc7fb,64'hb9ef9b20a887a698,64'h047dbe1bdc5c2e14,64'h15ba25eb47d1970b,
64'h064d2b36b592b1ba,64'hd9341d15b7db490e,64'hcf7500d8f76a5efe,64'h5e4bb2b1aa63a064,
64'hbdd7169e7c771904,64'h2474a3e4bb82a9d5,64'h2b1953f51993352f,64'h0000000080000000,
64'hf2a78e2633d89d74,64'h306a9ebec2d37535,64'h078cdff28fdeba24,64'h5732a953e12fd009,
64'h03019f8c5ffac78d,64'hc70965f0fe591a2e,64'ha2a2a91d423f5479,64'hae5253591bde074f,
64'h776fda6ab26dd0fc,64'hd7c1a5d80051efcd,64'h6ffa4109f2a940ca,64'h361d6230e328294a,
64'h677f2d42e7ac6c1b,64'ha8f89023d489f0e1,64'h4ae47916fec27627,64'h832a594f9e909747,
64'h88b38404fa95e091,64'hf692db7d4678e118,64'h02f367e3ad661c1a,64'hc24d5fc5fa01328c,
64'h67e541ea595d32db,64'hcc884007e2f06de6,64'h809a741e24309bc4,64'hcc72fe59d2b187bd,
64'hb7ebb438cc52b8ec,64'h896ffb80c6e620cb,64'h21303ba146df3c13,64'h632f689cda166c11,
64'hafbd6a245d1c6935,64'h3b93bb1b67ad75d1,64'h3be104974943ea75,64'hfefffffeffffff01,
64'h62ede5c3198e1ab5,64'h2903ed771a38edb8,64'hd84570bbe0daeca1,64'hb72f4c5e29bbab91,
64'hdcc9212aed37d080,64'hcea99570e08dd4d0,64'h42df2cbf4b4a18ce,64'h087a3bee02a7546f,
64'h054e3bba4d981250,64'hf22f71244084394c,64'h3dbc4c1c25dc4c9d,64'hee20087be15544ff,
64'hd239ddfd739c428c,64'hcae6bbab3a4fe778,64'h5658ff8b64b74cf5,64'h80eb1717fd252776,
64'h20ba8e254c483b13,64'hf5481698ba73fb2b,64'h04d780f218fdeb75,64'h74ec79564c5ff6cc,
64'he4e33045c5e63fd2,64'hcf7cd90a443d34bb,64'h23edf0dee2e170a0,64'hadd12f5a3e8cb858,
64'h326959b5ac958dd0,64'hc9a0e8b3beda486a,64'h7ba806cdbb52f7ea,64'hf25d958f531d031e,
64'heeb8b4f8e3b8c81b,64'h23a51f26dc154ea7,64'h58ca9fa9cc99a977,64'h0000000400000000,
64'h953c71389ec4eb99,64'h8354f5f7169ba9a7,64'h3c66ff947ef5d120,64'hb9954aa1097e8046,
64'h180cfc62ffd63c68,64'h384b2f8df2c8d16a,64'h151548ef11faa3c3,64'h72929acddef03a73,
64'hbb7ed358936e87dd,64'hbe0d2ec6028f7e62,64'h7fd20852954a064d,64'hb0eb118819414a4f,
64'h3bf96a1a3d6360d5,64'h47c48123a44f8703,64'h5723c8b9f613b136,64'h1952ca80f484ba34,
64'h459c202bd4af0484,64'hb496dbf133c708b9,64'h179b3f1d6b30e0d0,64'h126afe35d009945a,
64'h3f2a0f55cae996d5,64'h6442004517836f2a,64'h04d3a0f52184de1c,64'h6397f2d4958c3de2,
64'hbf5da1cb6295c75b,64'h4b7fdc0a37310654,64'h0981dd0b36f9e097,64'h197b44e9d0b36085,
64'h7deb5127e8e349a3,64'hdc9dd8dc3d6bae87,64'hdf0824bb4a1f53a7,64'hf7fffffefffff801,
64'h176f2e1bcc70d5a5,64'h481f6bb9d1c76dbf,64'hc22b85e506d76502,64'hb97a62f64ddd5c83,
64'he649095d69be83fa,64'h754cab8d046ea67a,64'h16f965fc5a50c66e,64'h43d1df70153aa378,
64'h2a71ddd26cc09280,64'h917b89290421ca59,64'hede260e22ee264e7,64'h710043e60aaa27f1,
64'h91ceeff19ce2145a,64'h5735dd5fd27f3bba,64'hb2c7fc5d25ba67a6,64'h0758b8c3e9293bac,
64'h05d4712b6241d897,64'haa40b4ccd39fd951,64'h26bc0790c7ef5ba8,64'ha763cab562ffb65d,
64'h271982352f31fe89,64'h7be6c85821e9a5d2,64'h1f6f86f8170b84ff,64'h6e897ad6f465c2bb,
64'h934acdae64ac6e7f,64'h4d0745a3f6d2434a,64'hdd403670da97bf4d,64'h92ecac8198e818e9,
64'h75c5a7ce1dc640d1,64'h1d28f937e0aa7537,64'hc654fd5064cd4bb6,64'h0000002000000000,
64'ha9e389c8f6275cc4,64'h1aa7afbcb4dd4d34,64'he337fca4f7ae88ff,64'hccaa550d4bf4022b,
64'hc067e317feb1e340,64'hc2597c7096468b4f,64'ha8aa47788fd51e18,64'h9494d671f781d395,
64'hdbf69ac99b743ee3,64'hf0697635147bf30b,64'hfe904297aa503265,64'h87588c45ca0a5273,
64'hdfcb50d2eb1b06a7,64'h3e24091f227c3816,64'hb91e45d1b09d89ae,64'hca965407a425d1a0,
64'h2ce10160a578241e,64'ha4b6df8e9e3845c3,64'hbcd9f8eb59870680,64'h9357f1ae804ca2d0,
64'hf9507aaf574cb6a7,64'h2210022bbc1b794d,64'h269d07a90c26f0e0,64'h1cbf96a7ac61ef0d,
64'hfaed0e6014ae3ad3,64'h5bfee053b988329e,64'h4c0ee859b7cf04b8,64'hcbda274e859b0428,
64'hef5a8942471a4d15,64'he4eec6e7eb5d7432,64'hf84125e050fa9d32,64'hbffffffeffffc001,
64'hbb7970de6386ad28,64'h40fb5dd08e3b6df6,64'h115c2f2e36bb280a,64'hcbd317b76eeae413,
64'h32484af24df41fc9,64'haa655c6b237533cd,64'hb7cb2fe2d2863370,64'h1e8efb82a9d51bbe,
64'h538eee94660493ff,64'h8bdc494c210e52c4,64'h6f13071877132731,64'h88021f3355513f85,
64'h8e777f90e710a2cc,64'hb9aeeb0093f9ddce,64'h963fe2ee2dd33d2b,64'h3ac5c61f4949dd60,
64'h2ea3895b120ec4b8,64'h5205a66b9cfeca83,64'h35e03c873f7add3f,64'h3b1e55b017fdb2e3,
64'h38cc11aa798ff447,64'hdf3642c40f4d2e8d,64'hfb7c37c0b85c27f8,64'h744bd6baa32e15d5,
64'h9a566d77256373f4,64'h683a2d21b6921a4e,64'hea01b38cd4bdfa62,64'h97656410c740c744,
64'hae2d3e73ee320685,64'he947c9bf0553a9b8,64'h32a7ea89266a5daa,64'h0000010000000000,
64'h4f1c4e4cb13ae61b,64'hd53d7de5a6ea69a0,64'h19bfe52ebd7447f1,64'h6552a8705fa01152,
64'h033f18c5f58f19fa,64'h12cbe38ab2345a72,64'h45523bc97ea8f0bb,64'ha4a6b393bc0e9ca4,
64'hdfb4d652dba1f712,64'h834bb1afa3df9851,64'hf48214c452819321,64'h3ac4623250529394,
64'hfe5a869d58d83532,64'hf12048fa13e1c0af,64'hc8f22e9284ec4d6b,64'h54b2a043212e8cfa,
64'h67080b062bc120ef,64'h25b6fc79f1c22e13,64'he6cfc75fcc3833fb,64'h9abf8d780265167c,
64'hca83d581ba65b531,64'h1080115ee0dbca67,64'h34e83d49613786ff,64'he5fcb53d630f7868,
64'hd7687307a571d691,64'hdff7029fcc4194ee,64'h607742cfbe7825be,64'h5ed13a7a2cd8213a,
64'h7ad44a1938d268a1,64'h277637465aeba189,64'hc2092f0987d4e989,64'hfffffffcfffe0003,
64'hdbcb86f81c35693b,64'h07daee8671db6fae,64'h8ae17971b5d94050,64'h5e98bdc177572092,
64'h924257936fa0fe47,64'h532ae35e1ba99e63,64'hbe597f1b94319b7b,64'hf477dc154ea8ddf0,
64'h9c7774a530249ff6,64'h5ee24a650872961c,64'h789838c6b8993985,64'h4010f99eaa89fc24,
64'h73bbfc8b3885165c,64'hcd7758099fceee6b,64'hb1ff17756e99e954,64'hd62e30fb4a4eeaff,
64'h751c4ad9907625bf,64'h902d335ee7f65416,64'haf01e43afbd6e9f7,64'hd8f2ad81bfed9717,
64'hc6608d54cc7fa237,64'hf9b216267a697462,64'hdbe1be0cc2e13fb9,64'ha25eb5d81970aea5,
64'hd2b36bbd2b1b9f9c,64'h41d16910b490d26d,64'h500d9c6da5efd309,64'hbb2b208a3a063a1c,
64'h7169f3a471903423,64'h4a3e4dff2a9d4db9,64'h953f544a3352ed4f,64'h0000080000000000,
64'h78e2726789d730d6,64'ha9ebef3337534cfa,64'hcdff2975eba23f88,64'h2a954385fd008a8d,
64'h19f8c62fac78cfd0,64'h965f1c5591a2d390,64'h2a91de4df54785d6,64'h25359ca2e074e51b,
64'hfda6b29cdd0fb88a,64'h1a5d8d811efcc284,64'ha410a629940c9901,64'hd623119382949c9f,
64'hf2d434f1c6c1a989,64'h890247d79f0e0571,64'h4791749a27626b52,64'ha595021b097467ce,
64'h384058345e090775,64'h2db7e3d08e117097,64'h367e3b0561c19fd1,64'hd5fc6bc41328b3dc,
64'h541eac13d32da982,64'h84008af706de5338,64'ha741ea4c09bc37f7,64'h2fe5a9f2187bc339,
64'hbb4398432b8eb482,64'hffb81504620ca76a,64'h03ba1680f3c12ded,64'hf689d3d366c109ce,
64'hd6a250ccc6934505,64'h3bb1ba33d75d0c47,64'h104978523ea74c42,64'hffffffeefff00011,
64'hde5c37c6e1ab49d2,64'h3ed774338edb7d70,64'h570bcb91aeca027c,64'hf4c5ee0dbab9048e,
64'h9212bc9f7d07f234,64'h99571af2dd4cf316,64'hf2cbf8e1a18cdbd3,64'ha3bee0b17546ef79,
64'he3bba52d8124ffac,64'hf712532a4394b0de,64'hc4c1c638c4c9cc25,64'h0087ccf7544fe11e,
64'h9ddfe45cc428b2dd,64'h6bbac052fe777352,64'h8ff8bbb074cf4a9b,64'hb17187e0527757f2,
64'ha8e256cf83b12df5,64'h81699afb3fb2a0ac,64'h780f21dcdeb74fb3,64'hc7956c13ff6cb8b2,
64'h33046aac63fd11b2,64'hcd90b13ad34ba309,64'hdf0df06c1709fdc2,64'h12f5aec5cb857523,
64'h959b5def58dcfcda,64'h0e8b4887a4869366,64'h806ce36f2f7e9846,64'hd9590456d031d0db,
64'h8b4f9d268c81a115,64'h51f26ffb54ea6dc6,64'ha9faa2559a976a74,64'h0000400000000000,
64'hc713933f4eb986ad,64'h4f5f799eba9a67cb,64'h6ff94bb55d11fc3a,64'h54aa1c30e8045467,
64'hcfc6317d63c67e80,64'hb2f8e2b08d169c7c,64'h548ef270aa3c2eaf,64'h29ace51803a728d7,
64'hed3594ede87dc449,64'hd2ec6c08f7e61420,64'h20853151a064c803,64'hb1188ca214a4e4f2,
64'h96a1a795360d4c41,64'h48123ec0f8702b84,64'h3c8ba4d33b135a8e,64'h2ca810dd4ba33e6b,
64'hc202c1a3f0483ba7,64'h6dbf1e85708b84b7,64'hb3f1d82c0e0cfe87,64'hafe35e2699459eda,
64'ha0f560a0996d4c0e,64'h200457bc36f299bc,64'h3a0f52654de1bfb3,64'h7f2d4f91c3de19c7,
64'hda1cc21e5c75a40b,64'hfdc0a82a10653b49,64'h1dd0b4079e096f68,64'hb44e9ea236084e69,
64'hb512866c349a2822,64'hdd8dd19fbae86237,64'h824bc291f53a6210,64'hffffff7eff800081,
64'hf2e1be3d0d5a4e8a,64'hf6bba19d76dbeb7f,64'hb85e5c8f765013de,64'ha62f7074d5c82469,
64'h9095e4ffe83f919c,64'hcab8d79aea6798ac,64'h965fc7140c66de91,64'h1df70590aa377bc3,
64'h1ddd29730927fd59,64'hb89299591ca586e9,64'h260e31cc264e6122,64'h043e67baa27f08f0,
64'heeff22ea214596e4,64'h5dd6029af3bb9a8d,64'h7fc5dd87a67a54d4,64'h8b8c3f0793babf8b,
64'h4712b6811d896fa3,64'h0b4cd7ddfd95055c,64'hc0790ee9f5ba7d95,64'h3cab60a5fb65c58a,
64'h982355641fe88d8f,64'h6c8589dc9a5d1842,64'hf86f8366b84fee0a,64'h97ad762e5c2ba918,
64'hacdaef7ec6e7e6cc,64'h745a443d24349b30,64'h03671b7d7bf4c22c,64'hcac822bc818e86d2,
64'h5a7ce938640d08a4,64'h8f937fdca7536e2e,64'h4fd512b1d4bb539b,64'h0002000000000000,
64'h389c9a0075cc3562,64'h7afbccf7d4d33e56,64'h7fca5dade88fe1cd,64'ha550e1894022a336,
64'h7e318bf11e33f3fa,64'h97c7158968b4e3db,64'ha477938751e17576,64'h4d6728c11d3946b7,
64'h69aca77643ee2241,64'h9763604dbf30a0fa,64'h04298a8e03264017,64'h88c46515a527278b,
64'hb50d3cadb06a6204,64'h4091f609c3815c1e,64'he45d269ad89ad46f,64'h654086eb5d19f357,
64'h10160d258241dd32,64'h6df8f42e845c25b5,64'h9f8ec1657067f433,64'h7f1af139ca2cf6cb,
64'h07ab0509cb6a606b,64'h0022bde2b794cddf,64'hd07a932b6f0dfd97,64'hf96a7c911ef0ce35,
64'hd0e610f8e3ad2052,64'hee0541578329da41,64'hee85a03cf04b7b40,64'ha274f516b0427343,
64'ha8943366a4d1410b,64'hec6e8d03d74311b2,64'h125e1493a9d3107c,64'hfffffbfefc000401,
64'h970df1ef6ad27449,64'hb5dd0cf2b6df5bf1,64'hc2f2e480b2809eeb,64'h317b83abae412343,
64'h84af280341fc8cdc,64'h55c6bcdd533cc55a,64'hb2fe38a46336f484,64'hefb82c8551bbde18,
64'heee94b98493feac8,64'hc494cacde52c3743,64'h30718e623273090f,64'h21f33dd513f84780,
64'h77f917580a2cb719,64'heeb014d99ddcd466,64'hfe2eec4033d2a69d,64'h5c61f8409dd5fc54,
64'h3895b40aec4b7d16,64'h5a66beefeca82ae0,64'h03c87755add3eca2,64'he55b0530db2e2c4f,
64'hc11aab24ff446c74,64'h642c4ee7d2e8c20d,64'hc37c1b3cc27f7049,64'hbd6bb176e15d48bc,
64'h66d77bfb373f365b,64'ha2d221ec21a4d97d,64'h1b38dbebdfa61160,64'h564115ea0c74368a,
64'hd3e749c52068451e,64'h7c9bfee93a9b716c,64'h7ea89590a5da9cd6,64'h0010000000000000,
64'hc4e4d004ae61ab0f,64'hd7de67c1a699f2ad,64'hfe52ed72447f0e65,64'h2a870c4f011519ab,
64'hf18c5f8bf19f9fcd,64'hbe38ac4f45a71ed4,64'h23bc9c3f8f0babab,64'h6b39460ae9ca35b6,
64'h4d653bb51f711205,64'hbb1b0271f98507cc,64'h214c5470193200b8,64'h462328b129393c54,
64'ha869e5728353101b,64'h048fb0501c0ae0ee,64'h22e934ddc4d6a371,64'h2a04375de8cf9ab5,
64'h80b0692c120ee990,64'h6fc7a17722e12da5,64'hfc760b2f833fa194,64'hf8d789d15167b655,
64'h3d58284e5b530358,64'h0115ef15bca66ef8,64'h83d49961786fecb2,64'hcb53e48ff78671a1,
64'h873087cd1d69028a,64'h702a0ac3194ed201,64'h742d01ee825bd9f9,64'h13a7a8ba82139a13,
64'h44a19b3a268a0853,64'h63746825ba188d89,64'h92f0a49d4e9883e0,64'hffffdffee0002001,
64'hb86f8f7f5693a244,64'haee8679ab6fadf83,64'h1797240b9404f752,64'h8bdc1d5e72091a17,
64'h2579401e0fe466dc,64'hae35e6ec99e62ace,64'h97f1c52819b7a41b,64'h7dc164318ddef0b9,
64'h774a5cc949ff5639,64'h24a656752961ba12,64'h838c731293984877,64'h0f99eea99fc23bff,
64'hbfc8bac35165b8c5,64'h7580a6d3eee6a329,64'hf17762089e9534e1,64'he30fc206eeafe29e,
64'hc4ada058625be8af,64'hd335f781654156fe,64'h1e43baad6e9f6510,64'h2ad8298dd9716271,
64'h08d5592dfa23639a,64'h2162774197461065,64'h1be0d9ec13fb8242,64'heb5d8bbc0aea45db,
64'h36bbdfdcb9f9b2d5,64'h16910f660d26cbe3,64'hd9c6df5efd308b00,64'hb208af5263a1b44e,
64'h9f3a4e2f034228ea,64'he4dff74cd4db8b5d,64'hf544ac882ed4e6ad,64'h0080000000000000,
64'h2726802b730d5872,64'hbef33e1334cf9562,64'hf2976b9923f87321,64'h5438627908a8cd57,
64'h8c62fc668cfcfe61,64'hf1c5627f2d38f69b,64'h1de4e1fd785d5d57,64'h59ca305a4e51adad,
64'h6b29ddaafb889026,64'hd8d81394cc283e5b,64'h0a62a381c99005bf,64'h3119458b49c9e29e,
64'h434f2b991a9880d3,64'h247d8280e0570770,64'h1749a6ef26b51b87,64'h5021baf0467cd5a7,
64'h0583496490774c7c,64'h7e3d0bbc17096d25,64'he3b0598319fd0c99,64'hc6bc4e918b3db2a1,
64'heac14273da981abf,64'h08af78ade53377c0,64'h1ea4cb0fc37f658c,64'h5a9f2485bc338d02,
64'h39843e6ceb48144c,64'h8150561bca769005,64'ha1680f7712decfc5,64'h9d3d45d4109cd098,
64'h250cd9d334504296,64'h1ba34130d0c46c45,64'h978524ee74c41efc,64'hfffefffe00010001,
64'hc37c7bffb49d121b,64'h77433cdab7d6fc13,64'hbcb9205ca027ba90,64'h5ee0eaf79048d0b4,
64'h2bca00f17f2336df,64'h71af3769cf31566b,64'hbf8e2944cdbd20d4,64'hee0b218f6ef785c5,
64'hba52e64d4ffab1c5,64'h2532b3aa4b0dd08f,64'h1c6398989cc243b4,64'h7ccf754cfe11dff8,
64'hfe45d61f8b2dc623,64'hac0536a277351945,64'h8bbb104bf4a9a701,64'h187e103e757f14e9,
64'h256d02c912df4572,64'h99afbc112a0ab7ea,64'hf21dd56b74fb2880,64'h56c14c6fcb8b1387,
64'h46aac96fd11b1cd0,64'h0b13ba0dba308327,64'hdf06cf609fdc1210,64'h5aec5de757522ed1,
64'hb5defee6cfcd96a7,64'hb4887b3069365f18,64'hce36fafde98457fa,64'h90457a981d0da26b,
64'hf9d2717c1a11474c,64'h26ffba6da6dc5ae1,64'haa25644876a73561,64'h0400000000000000,
64'h3934015c986ac38f,64'hf799f09ea67cab0b,64'h94bb5cd01fc39901,64'ha1c313ca45466ab6,
64'h6317e33867e7f304,64'h8e2b140069c7b4d1,64'hef270febc2eaeab8,64'hce5182d4728d6d66,
64'h594eed5adc44812d,64'hc6c09cac6141f2d2,64'h53151c0e4c802df8,64'h88ca2c5b4e4f14ef,
64'h1a795ccad4c40696,64'h23ec140802b83b7f,64'hba4d377935a8dc38,64'h810dd78433e6ad36,
64'h2c1a4b2483ba63e0,64'hf1e85de3b84b6925,64'h1d82cc1fcfe864c1,64'h35e2749259ed9502,
64'h560a13a5d4c0d5f1,64'h457bc56f299bbe00,64'hf526587e1bfb2c60,64'hd4f9242fe19c680e,
64'hcc21f3685a40a25f,64'h0a82b0e253b48024,64'h0b407bbd96f67e23,64'he9ea2ea484e684bc,
64'h2866ce9aa28214af,64'hdd1a098686236228,64'hbc292777a620f7dc,64'hfff7fff700080001,
64'h1be3e003a4e890d2,64'hba19e6d8beb7e095,64'he5c902ea013dd47b,64'hf70757be8246859e,
64'h5e50078cf919b6f7,64'h8d79bb51798ab355,64'hfc714a2b6de9069b,64'h70590c8277bc2e21,
64'hd297326f7fd58e23,64'h29959d53586e8477,64'he31cc4c4e6121da0,64'he67baa6af08effbd,
64'hf22eb103596e3111,64'h6029b518b9a8ca23,64'h5dd88263a54d3804,64'hc3f081f3abf8a748,
64'h2b68164996fa2b8f,64'hcd7de08d5055bf4c,64'h90eeab62a7d943f9,64'hb60a63805c589c36,
64'h35564b8088d8e67e,64'h589dd06dd1841938,64'hf8367b0afee0907a,64'hd762ef3cba917686,
64'haef7f73b7e6cb533,64'ha443d98849b2f8bb,64'h71b7d7f54c22bfca,64'h822bd4c4e86d1354,
64'hce938be7d08a3a59,64'h37fdd36e36e2d707,64'h512b2248b539ab03,64'h2000000000000000,
64'hc9a00ae5c3561c77,64'hbccf84fc33e55851,64'ha5dae684fe1cc804,64'h0e189e572a3355ab,
64'h18bf19c63f3f981d,64'h7158a0074e3da684,64'h79387f65175755b9,64'h728c16a9946b6b2a,
64'hca776ad8e2240966,64'h3604e5690a0f968a,64'h98a8e07464016fbe,64'h465162de7278a774,
64'hd3cae656a62034b0,64'h1f60a04115c1dbf7,64'hd269bbcead46e1bb,64'h086ebc259f3569ac,
64'h60d259251dd31eff,64'h8f42ef24c25b4921,64'hec1660fe7f432608,64'haf13a493cf6ca80f,
64'hb0509d30a606af86,64'h2bde2b7b4cddeffe,64'ha932c3f7dfd962f9,64'ha7c921850ce3406a,
64'h610f9b48d20512f2,64'h541587129da40120,64'h5a03ddecb7b3f118,64'h4f51752b273425d9,
64'h433674d61410a577,64'he8d04c3a311b113a,64'he1493bc23107bedb,64'hffbfffbf00400001,
64'hdf1f001d27448690,64'hd0cf36caf5bf04a3,64'h2e48175709eea3d1,64'hb83abdfb12342ce9,
64'hf2803c69c8cdb7b6,64'h6bcdda8fcc559aa4,64'he38a51626f4834d1,64'h82c86416bde17105,
64'h94b99381feac7112,64'h4cacea9bc37423b7,64'h18e6262e3090ecf9,64'h33dd535e8477fde1,
64'h91758821cb718881,64'h014da8c8cd465115,64'heec4131f2a69c01e,64'h1f840fa35fc53a3a,
64'h5b40b24db7d15c77,64'h6bef047082adfa5a,64'h87755b193eca1fc4,64'hb0531c07e2c4e1ab,
64'haab25c0546c733ef,64'hc4ee83708c20c9be,64'hc1b3d85ef70483c9,64'hbb1779ebd48bb42a,
64'h77bfb9e0f365a993,64'h221ecc474d97c5d3,64'h8dbebfad6115fe4d,64'h115ea62b43689a9c,
64'h749c5f448451d2c2,64'hbfee9b72b716b837,64'h89591247a9cd5816,64'h00000000ffffffff,
64'h4d0057341ab0e3b2,64'he67c27e69f2ac283,64'h2ed7342cf0e6401b,64'h70c4f2b9519aad58,
64'hc5f8ce31f9fcc0e8,64'h8ac5003d71ed341d,64'hc9c3fb2bbabaadc5,64'h9460b54fa35b594d,
64'h53bb56cd11204b2a,64'hb0272b49507cb44f,64'hc54703a7200b7dec,64'h328b16f593c53b9e,
64'h9e5732bb3101a57a,64'hfb050208ae0edfb8,64'h934dde7b6a370dd2,64'h4375e12cf9ab4d60,
64'h0692c92bee98f7f5,64'h7a17792a12da4904,64'h60b307fafa193039,64'h789d24a37b654073,
64'h8284e98a30357c2b,64'h5ef15bdb66ef7fef,64'h49961fc3fecb17c3,64'h3e490c2d671a034b,
64'h087cda499028978d,64'ha0ac3896ed2008fe,64'hd01eef67bd9f88be,64'h7a8ba95b39a12ec6,
64'h19b3a6b2a0852bb6,64'h468261d888d889c9,64'h0a49de18883df6d1,64'hfdfffdff02000001,
64'hf8f800ef3a24347a,64'h8679b65dadf82512,64'h7240bab94f751e87,64'hc1d5efdd91a16743,
64'h9401e355466dbda9,64'h5e6ed48162acd51d,64'h1c528b1a7a41a681,64'h164320b9ef0b8824,
64'ha5cc9c13f563888c,64'h656754e01ba11db6,64'hc7313171848767c8,64'h9eea9af523bfef07,
64'h8bac41125b8c4404,64'h0a6d46466a3288a8,64'h76209900534e00e9,64'hfc207d1afe29d1d0,
64'hda05926fbe8ae3b6,64'h5f782387156fd2cd,64'h3baad8cdf650fe1c,64'h8298e04416270d53,
64'h5592e02f36399f73,64'h27741b8a61064dea,64'h0d9ec2fdb8241e42,64'hd8bbcf63a45da14b,
64'hbdfdcf0a9b2d4c95,64'h10f6623b6cbe2e97,64'h6df5fd6f08aff264,64'h8af5315a1b44d4e0,
64'ha4e2fa27228e960d,64'hff74db9ab8b5c1b3,64'h4ac892414e6ac0ac,64'h00000007fffffff8,
64'h6802b9a2d5871d8e,64'h33e13f3bf9561411,64'h76b9a168873200d7,64'h862795cd8cd56abd,
64'h2fc67195cfe6073a,64'h562801ef8f69a0e4,64'h4e1fd963d5d56e22,64'ha305aa811adaca64,
64'h9ddab66a8902594e,64'h81395a4f83e5a273,64'h2a381d3f005bef5a,64'h9458b7ad9e29dcef,
64'hf2b995dd880d2bcc,64'hd828104c7076fdb9,64'h9a6ef3df51b86e8c,64'h1baf0969cd5a6afe,
64'h3496495f74c7bfa8,64'hd0bbc95396d2481d,64'h05983fdad0c981c5,64'hc4e9251edb2a0395,
64'h14274c5581abe154,64'hf78adedd377bff76,64'h4cb0fe21f658be16,64'hf248616c38d01a57,
64'h43e6d24c8144bc68,64'h0561c4bc690047eb,64'h80f77b43ecfc45ea,64'hd45d4adccd09762d,
64'hcd9d359504295db0,64'h34130ec646c44e46,64'h524ef0c441efb688,64'hefffefff10000001,
64'hc7c00780d121a3c9,64'h33cdb2f16fc1288c,64'h9205d5cd7ba8f435,64'h0eaf7ef28d0b3a12,
64'ha00f1aae336ded44,64'hf376a40d1566a8e6,64'he29458d3d20d3408,64'hb21905cf785c4120,
64'h2e64e0a4ab1c445b,64'h2b3aa703dd08edad,64'h39898b92243b3e3a,64'hf754d7ad1dff7834,
64'h5d620896dc62201c,64'h536a323351944540,64'hb104c8059a700745,64'he103e8def14e8e79,
64'hd02c9383f4571daa,64'hfbc11c3aab7e9666,64'hdd56c670b287f0df,64'h14c70224b1386a94,
64'hac97017bb1ccfb96,64'h3ba0dc5408326f4f,64'h6cf617edc120f210,64'hc5de7b2322ed0a52,
64'hefee7859d96a64a3,64'h87b311db65f174b8,64'h6fafeb7b457f931d,64'h57a98ad4da26a6fc,
64'h2717d13e1474b063,64'hfba6dcdcc5ae0d91,64'h5644920c7356055e,64'h0000003fffffffc0,
64'h4015cd19ac38ec6d,64'h9f09f9e0cab0a087,64'hb5cd0b47399006b5,64'h313cae7066ab55e4,
64'h7e338caf7f3039cf,64'hb1400f7e7b4d071e,64'h70fecb20aeab710e,64'h182d540dd6d6531b,
64'heed5b3584812ca6c,64'h09cad2801f2d1394,64'h51c0e9f902df7acf,64'ha2c5bd70f14ee774,
64'h95ccaef340695e59,64'hc140826983b7edc2,64'hd3779efe8dc3745c,64'hdd784b4e6ad357f0,
64'ha4b24afca63dfd3f,64'h85de4aa2b69240e2,64'h2cc1fed6864c0e28,64'h274928fcd9501ca2,
64'ha13a62ac0d5f0aa0,64'hbc56f6f0bbdffba9,64'h6587f111b2c5f0ae,64'h92430b68c680d2b1,
64'h1f3692660a25e33e,64'h2b0e25e348023f58,64'h07bbda2367e22f4c,64'ha2ea56ec684bb162,
64'h6ce9acae214aed7a,64'ha09876333622722f,64'h927786240f7db43e,64'h7fff7fff80000001,
64'h3e003c0c890d1e42,64'h9e6d978c7e09445f,64'h902eae6fdd47a1a4,64'h757bf7946859d090,
64'h0078d5769b6f6a1b,64'h9bb5206fab354729,64'h14a2c6a59069a039,64'h90c82e80c2e208fb,
64'h7327052658e222d7,64'h59d5381fe8476d67,64'hcc4c5c9221d9f1cf,64'hbaa6bd6feffbc199,
64'heb1044b8e31100de,64'h9b51919c8ca229fe,64'h88264031d3803a23,64'h081f46fe8a7473c1,
64'h81649c25a2b8ed4a,64'hde08e1dc5bf4b329,64'heab6338b943f86f2,64'ha638112589c354a0,
64'h64b80be28e67dcab,64'hdd06e2a141937a77,64'h67b0bf710907907d,64'h2ef3d91f1768528a,
64'h7f73c2d5cb532511,64'h3d988edf2f8ba5bc,64'h7d7f5bdd2bfc98e5,64'hbd4c56a8d13537de,
64'h38be89f1a3a58317,64'hdd36e6ed2d706c81,64'hb22490659ab02aee,64'h000001fffffffe00,
64'h00ae68cf61c76366,64'hf84fcf0a55850434,64'hae685a3ecc8035a3,64'h89e57384355aaf1f,
64'hf19c657ef981ce75,64'h8a007bf8da6838eb,64'h87f65908755b886d,64'hc16aa06eb6b298d8,
64'h76ad9ac940965359,64'h4e569400f9689ca0,64'h8e074fca16fbd676,64'h162deb8c8a773b9b,
64'hae65779e034af2c4,64'h0a0413521dbf6e0a,64'h9bbcf7fa6e1ba2da,64'hebc25a79569abf7a,
64'h259257ea31efe9f3,64'h2ef25519b492070c,64'h660ff6b53260713f,64'h3a4947e7ca80e50f,
64'h09d315656af854fb,64'he2b7b78adeffdd43,64'h2c3f8890962f856d,64'h92185b4a34069584,
64'hf9b49330512f19f0,64'h58712f1b4011fabf,64'h3dded11b3f117a60,64'h1752b768425d8b0b,
64'h674d65740a576bcd,64'h04c3b19eb1139173,64'h93bc31247beda1ec,64'hfffbffff00000005,
64'hf001e0654868f20f,64'hf36cbc67f04a22f4,64'h81757382ea3d0d1c,64'habdfbca642ce847d,
64'h03c6abb4db7b50d8,64'hdda9038159aa3944,64'ha516352c834d01c8,64'h8641740a171047d4,
64'h99382935c71116b5,64'hcea9c101423b6b36,64'h6262e4970ecf8e72,64'hd535eb847fde0cc3,
64'h588225ce188806e9,64'hda8c8ce865114fec,64'h413201929c01d114,64'h40fa37f453a39e08,
64'h0b24e13115c76a4c,64'hf0470ee8dfa59942,64'h55b19c63a1fc3789,64'h31c089314e1aa4fb,
64'h25c05f17733ee555,64'he83715100c9bd3b2,64'h3d85fb8b483c83e5,64'h779ec8f9bb42944f,
64'hfb9e16b15a992885,64'hecc476fa7c5d2ddf,64'hebfadeec5fe4c725,64'hea62b54b89a9beeb,
64'hc5f44f8e1d2c18b7,64'he9b7376f6b836402,64'h91248331d581576b,64'h00000ffffffff000,
64'h0573467b0e3b1b30,64'hc27e7859ac282199,64'h7342d1fb6401ad13,64'h4f2b9c25aad578f4,
64'h8ce32bfecc0e73a1,64'h5003dfcad341c754,64'h3fb2c847aadc4364,64'h0b55037bb594c6ba,
64'hb56cd64d04b29ac5,64'h72b4a009cb44e4fe,64'h703a7e54b7deb3ac,64'hb16f5c6453b9dcd8,
64'h732bbcf51a57961b,64'h50209a90edfb7050,64'hdde7bfd770dd16cc,64'h5e12d3d1b4d5fbc9,
64'h2c92bf528f7f4f97,64'h7792a8cea490385f,64'h307fb5ac930389f5,64'hd24a3f3f54072877,
64'h4e98ab2b57c2a7d8,64'h15bdbc5df7feea11,64'h61fc4485b17c2b67,64'h90c2da55a034ac1c,
64'hcda499898978cf79,64'hc38978dc008fd5f6,64'heef688daf88bd2ff,64'hba95bb4212ec5858,
64'h3a6b2ba352bb5e65,64'h261d8cf5889c8b98,64'h9de18927df6d0f5c,64'hffdfffff00000021,
64'h800f033143479071,64'h9b65e34682511799,64'h0bab9c1b51e868dc,64'h5efde537167423e3,
64'h1e355da6dbda86c0,64'hed481c10cd51ca1a,64'h28b1a9691a680e3b,64'h320ba054b8823e9c,
64'hc9c149b23888b5a4,64'h754e081011db59aa,64'h131724bb767c738d,64'ha9af5c29fef06612,
64'hc4112e72c4403746,64'hd4646749288a7f5a,64'h09900c96e00e889e,64'h07d1bfa49d1cf03e,
64'h59270988ae3b5260,64'h8238774dfd2cca09,64'had8ce31f0fe1bc46,64'h8e04498b70d527d7,
64'h2e02f8bc99f72aa7,64'h41b8a88764de9d89,64'hec2fdc5b41e41f27,64'hbcf647d0da14a275,
64'hdcf0b591d4c94421,64'h6623b7dae2e96ef1,64'h5fd6f769ff263921,64'h5315aa634d4df751,
64'h2fa27c76e960c5b2,64'h4db9bb825c1b2009,64'h89241992ac0abb54,64'h00007fffffff8000,
64'h2b9a33d871d8d980,64'h13f3c2d361410cc2,64'h9a168fde200d6895,64'h795ce12f56abc79e,
64'h67195ffa60739d04,64'h801efe589a0e3a9e,64'hfd96423e56e21b1f,64'h5aa81bddaca635d0,
64'hab66b26d2594d623,64'h95a500515a2727ed,64'h81d3f2a8bef59d5d,64'h8b7ae3279dcee6bb,
64'h995de7abd2bcb0d5,64'h8104d4896fdb827e,64'hef3dfec186e8b65a,64'hf0969e8fa6afde46,
64'h6495fa957bfa7cb7,64'hbc9546782481c2f5,64'h83fdad65981c4fa7,64'h9251fa00a03943b2,
64'h74c5595cbe153ebe,64'hadede2efbff75088,64'h0fe224308be15b35,64'h8616d2b101a560dc,
64'h6d24cc524bc67bc2,64'h1c4bc6e6047eafaa,64'h77b446dec45e97f1,64'hd4adda159762c2bb,
64'hd3595d1b95daf327,64'h30ec67ad44e45cbf,64'hef0c4942fb687adc,64'hfeffffff00000101,
64'h0078198e1a3c8384,64'hdb2f1a381288bcc4,64'h5d5ce0da8f4346e0,64'hf7ef29bab3a11f16,
64'hf1aaed36ded43600,64'h6a40e08d6a8e50c9,64'h458d4b49d34071d7,64'h905d02a6c411f4df,
64'h4e0a4d97c445ad1a,64'haa7040838edacd4d,64'h98b925dbb3e39c68,64'h4d7ae154f783308b,
64'h2089739c2201ba2a,64'ha3233a4f4453faca,64'h4c8064b7007444f0,64'h3e8dfd24e8e781f0,
64'hc9384c4771da92fe,64'h11c3ba73e9665044,64'h6c6718fd7f0de22b,64'h70224c5f86a93eb4,
64'h7017c5e5cfb95537,64'h0dc5443d26f4ec46,64'h617ee2e10f20f931,64'he7b23e8bd0a513a3,
64'he785ac94a64a2102,64'h311dbeda174b7785,64'hfeb7bb51f931c906,64'h98ad531c6a6fba86,
64'h7d13e3b84b062d8f,64'h6dcddc14e0d90046,64'h4920cc996055da9c,64'h0003fffffffc0000,
64'h5cd19ec48ec6cbff,64'h9f9e169b0a086610,64'hd0b47ef5006b44a4,64'hcae7097db55e3ced,
64'h38caffd6039ce81d,64'h00f7f2c8d071d4ec,64'hecb211f9b710d8f1,64'hd540deef6531ae7e,
64'h5b35936e2ca6b113,64'had28028ed1393f64,64'h0e9f9549f7aceae4,64'h5bd71940ee7735d4,
64'hcaef3d6295e586a4,64'h0826a44f7edc13ec,64'h79eff6133745b2c9,64'h84b4f484357ef229,
64'h24afd4aedfd3e5b5,64'he4aa33c6240e17a3,64'h1fed6b30c0e27d34,64'h928fd00901ca1d8c,
64'ha62acae8f0a9f5ed,64'h6f6f1782ffba843b,64'h7f1121845f0ad9a8,64'h30b6958c0d2b06dc,
64'h692662955e33de0d,64'he25e373023f57d50,64'hbda236f922f4bf85,64'ha56ed0b2bb1615d2,
64'h9acae8e2aed79932,64'h87633d6b2722e5f7,64'h78624a1edb43d6d9,64'hf7ffffff00000801,
64'h03c0cc70d1e41c20,64'hd978d1c69445e61a,64'heae706d67a1a36fe,64'hbf794ddc9d08f8a9,
64'h8d5769bdf6a1aff9,64'h5207046e54728645,64'h2c6a5a509a038eb6,64'h82e8153a208fa6f4,
64'h70526cc0222d68ce,64'h5382042176d66a63,64'hc5c92ee19f1ce33c,64'h6bd70aa9bc198456,
64'h044b9ce2100dd14f,64'h1919d27f229fd64b,64'h640325ba03a2277e,64'hf46fe928473c0f7f,
64'h49c262418ed497ea,64'h8e1dd39f4b328220,64'h6338c7eef86f1155,64'h811262ff3549f59d,
64'h80be2f317dcaa9b5,64'h6e2a21e937a76230,64'h0bf7170b7907c985,64'h3d91f46585289d11,
64'h3c2d64ac32510809,64'h88edf6d1ba5bbc27,64'hf5bdda96c98e4829,64'hc56a98e7537dd42c,
64'he89f1dc558316c75,64'h6e6ee0aa06c8022d,64'h490664cd02aed4de,64'h001fffffffe00000,
64'he68cf62676365ff6,64'hfcf0b4dc5043307c,64'h85a3f7ae035a251a,64'h57384bf3aaf1e762,
64'hc657feb11ce740e7,64'h07bf9646838ea760,64'h65908fd4b886c781,64'haa06f781298d73ea,
64'hd9ac9b7365358896,64'h6940147b89c9fb1b,64'h74fcaa4fbd675720,64'hdeb8ca0973b9ae9e,
64'h5779eb1aaf2c351a,64'h4135227bf6e09f60,64'hcf7fb09cba2d9645,64'h25a7a425abf79144,
64'h257ea577fe9f2da7,64'h25519e382070bd11,64'hff6b59860713e9a0,64'h947e804c0e50ec5c,
64'h3156574c854faf63,64'h7b78bc1afdd421d5,64'hf8890c25f856cd3d,64'h85b4ac61695836df,
64'h493314adf19ef065,64'h12f1b9881fabea79,64'hed11b7ce17a5fc23,64'h2b76859ad8b0ae8b,
64'hd657471976bcc98c,64'h3b19eb5d39172fb4,64'hc31250f9da1eb6c5,64'hbfffffff00004001,
64'h1e0663868f20e100,64'hcbc68e3aa22f30ca,64'h573836bad0d1b7e9,64'hfbca6ee9e847c543,
64'h6abb4df3b50d7fc4,64'h90382374a3943226,64'h6352d285d01c75af,64'h1740a9d5047d379c,
64'h82936604116b466d,64'h9c10210db6b35316,64'h2e497712f8e719da,64'h5eb85550e0cc22ad,
64'h225ce710806e8a78,64'hc8ce93f914feb258,64'h20192dd31d113bed,64'ha37f494939e07bf1,
64'h4e13120e76a4bf4e,64'h70ee9cfe599410fc,64'h19c63f7ac3788aa5,64'h089317fdaa4face4,
64'h05f1798fee554da4,64'h71510f4cbd3b117d,64'h5fb8b85bc83e4c28,64'hec8fa32d2944e887,
64'he16b256292884047,64'h476fb691d2dde134,64'hadeed4bd4c724141,64'h2b54c7409beea15a,
64'h44f8ee31c18b63a1,64'h7377055336401165,64'h4833266a1576a6ee,64'h00ffffffff000000,
64'h3467b13ab1b2ffa9,64'he785a6e9821983d9,64'h2d1fbd741ad128cc,64'hb9c25f9f578f3b0e,
64'h32bff58ee73a0732,64'h3dfcb2341c753b00,64'h2c847ea8c4363c05,64'h5037bc0e4c6b9f4b,
64'hcd64dba129ac44aa,64'h4a00a3df4e4fd8d5,64'ha7e55280eb3ab8fd,64'hf5c650519dcd74ea,
64'hbbcf58d77961a8ce,64'h09a913e1b704fafe,64'h7bfd84ebd16cb222,64'h2d3d212e5fbc8a1f,
64'h2bf52bc0f4f96d37,64'h2a8cf1c20385e887,64'hfb5acc37389f4cf9,64'ha3f40264728762dc,
64'h8ab2ba652a7d7b17,64'hdbc5e0daeea10ea5,64'hc4486136c2b669e1,64'h2da5630f4ac1b6f4,
64'h4998a5718cf78326,64'h978dcc40fd5f53c8,64'h688dbe77bd2fe111,64'h5bb42cd7c5857457,
64'hb2ba38d1b5e64c5a,64'hd8cf5aeac8b97d9f,64'h189287d4d0f5b622,64'hfffffffd00020003,
64'hf0331c3479070800,64'h5e3471db1179864a,64'hb9c1b5d8868dbf46,64'hde537756423e2a11,
64'h55da6fa0a86bfe1d,64'h81c11ba91ca1912c,64'h1a96943180e3ad75,64'hba054ea823e9bce0,
64'h149b30248b5a3364,64'he0810871b59a98ac,64'h724bb898c738cecf,64'hf5c2aa8906611566,
64'h12e73885037453bf,64'h46749fcea7f592ba,64'h00c96e99e889df67,64'h1bfa4a4ecf03df83,
64'h70989075b525fa6e,64'h8774e7f5cca087dd,64'hce31fbd61bc45528,64'h4498bfed527d6720,
64'h2f8bcc7f72aa6d20,64'h8a887a68e9d88be5,64'hfdc5c2e041f2613e,64'h647d19704a274431,
64'h0b592b1b94420231,64'h3b7db49096ef099e,64'h6f76a5ef63920a03,64'h5aa63a05df750acf,
64'h27c771900c5b1d06,64'h9bb82a9cb2008b25,64'h41993352abb5376e,64'h07fffffff8000000,
64'ha33d89d68d97fd47,64'h3c2d375310cc1ec1,64'h68fdeba1d689465f,64'hce12fcffbc79d86b,
64'h95ffac7839d0398f,64'hefe591a1e3a9d7ff,64'h6423f54721b1e027,64'h81bde074635cfa56,
64'h6b26dd0f4d62254a,64'h50051efc727ec6a6,64'h3f2a940c59d5c7e3,64'hae328293ee6ba749,
64'hde7ac6c0cb0d466b,64'h4d489f0db827d7f0,64'hdfec27618b65910d,64'h69e90973fde450f7,
64'h5fa95e08a7cb69b7,64'h54678e111c2f4437,64'hdad661c0c4fa67c1,64'h1fa01328943b16db,
64'h5595d32d53ebd8b4,64'hde2f06dd75087522,64'h224309bc15b34f02,64'h6d2b187b560db79f,
64'h4cc52b8e67bc192e,64'hbc6e620beafa9e3c,64'h446df3c0e97f0885,64'hdda166c02c2ba2b6,
64'h95d1c692af3262cb,64'hc67ad75c45cbecf2,64'hc4943ea687adb110,64'hffffffef00100011,
64'h8198e1aac8383ff9,64'hf1a38eda8bcc324e,64'hce0daec9346dfa2b,64'hf29bbab811f15082,
64'haed37d07435ff0e6,64'h0e08dd4ce50c895c,64'hd4b4a18c071d6ba8,64'hd02a75461f4de6fb,
64'ha4d981245ad19b20,64'h04084394acd4c559,64'h925dc4c939c67675,64'hae15544f3308ab29,
64'h9739c4281ba29df8,64'h33a4fe773fac95ce,64'h064b74cf444efb38,64'hdfd25276781efc18,
64'h84c483b0a92fd36d,64'h3ba73fb265043ee4,64'h718fdeb6de22a93a,64'h24c5ff6c93eb38fe,
64'h7c5e63fc955368ff,64'h5443d34b4ec45f24,64'hee2e17090f9309e9,64'h23e8cb85513a2185,
64'h5ac958dca2101188,64'hdbeda485b7784cef,64'h7bb52f7e1c905015,64'hd531d030fba85676,
64'h3e3b8c8162d8e82f,64'hddc154e990045924,64'h0cc99a975da9bb6e,64'h3fffffffc0000000,
64'h19ec4eb96cbfea33,64'he169ba998660f607,64'h47ef5d11b44a32f5,64'h7097e803e3cec352,
64'haffd63c5ce81cc74,64'h7f2c8d161d4ebff1,64'h211faa3c0d8f0135,64'h0def03a71ae7d2ac,
64'h5936e87d6b112a4d,64'h8028f7e593f6352e,64'hf954a063ceae3f17,64'h719414a4735d3a43,
64'hf3d6360c586a3352,64'h6a44f86fc13ebf7e,64'hff613b125b2c8862,64'h4f484ba2ef2287b5,
64'hfd4af0473e5b4db6,64'ha33c708ae17a21b6,64'hd6b30e0c27d33e02,64'hfd009944a1d8b6d8,
64'hacae996c9f5ec59e,64'hf17836f1a843a90a,64'h12184de1ad9a780f,64'h6958c3ddb06dbcf5,
64'h66295c753de0c96e,64'he373106457d4f1db,64'h236f9e094bf84426,64'hed0b3607615d15aa,
64'hae8e349979931654,64'h33d6bae82e5f678a,64'h24a1f53a3d6d887a,64'hffffff7f00800081,
64'h0cc70d5a41c1ffc4,64'h8d1c76db5e619269,64'h706d764fa36fd152,64'h94ddd5c78f8a8409,
64'h769be83f1aff872b,64'h7046ea6728644ae0,64'ha5a50c6638eb5d3a,64'h8153aa36fa6f37d2,
64'h26cc0927d68cd8fb,64'h20421ca566a62ac8,64'h92ee264dce33b3a4,64'h70aaa27e98455943,
64'hb9ce2144dd14efbc,64'h9d27f3bafd64ae6f,64'h325ba67a2277d9c0,64'hfe9293b9c0f7e0ba,
64'h26241d89497e9b64,64'hdd39fd942821f71f,64'h8c7ef5b9f11549cd,64'h262ffb659f59c7ef,
64'he2f31fe7aa9b47f5,64'ha21e9a5c7622f91e,64'h7170b84f7c984f41,64'h1f465c2b89d10c27,
64'hd64ac6e710808c3e,64'hdf6d2433bbc26772,64'hdda97bf3e48280a5,64'ha98e818ddd42b3aa,
64'hf1dc640c16c74177,64'hee0aa7528022c91a,64'h664cd4baed4ddb70,64'hfffffffeffffffff,
64'hcf6275cb65ff5198,64'h0b4dd4d33307b031,64'h3f7ae88fa25197a6,64'h84bf40221e761a8d,
64'h7feb1e33740e639b,64'hf96468b3ea75ff85,64'h08fd51e16c7809a7,64'h6f781d38d73e9560,
64'hc9b743ed58895266,64'h0147bf309fb1a96c,64'hcaa503257571f8b1,64'h8ca0a5269ae9d215,
64'h9eb1b069c3519a89,64'h5227c38109f5fbed,64'hfb09d899d9644309,64'h7a425d1979143da6,
64'hea578240f2da6da9,64'h19e3845c0bd10dab,64'hb59870673e99f00a,64'he804ca2c0ec5b6b9,
64'h6574cb69faf62ceb,64'h8bc1b794421d4849,64'h90c26f0d6cd3c078,64'h4ac61ef0836de7a5,
64'h314ae3acef064b6d,64'h1b988329bea78ed1,64'h1b7cf04b5fc2212f,64'h6859b0420ae8ad49,
64'h7471a4d0cc98b29b,64'h9eb5d74272fb3c4f,64'h250fa9d2eb6c43cf,64'hfffffbff04000401,
64'h66386ad20e0ffe20,64'h68e3b6def30c9344,64'h836bb2801b7e8a8d,64'ha6eeae407c542044,
64'hb4df41fbd7fc3955,64'h8237533c432256fd,64'h2d286336c75ae9cb,64'h0a9d51bbd379be8c,
64'h3660493fb466c7d7,64'h0210e52c3531563f,64'h97713272719d9d1c,64'h855513f7c22aca15,
64'hce710a2be8a77ddb,64'he93f9ddbeb257374,64'h92dd33d213becdff,64'hf4949dd507bf05c9,
64'h3120ec4b4bf4db1f,64'he9cfeca7410fb8f2,64'h63f7add388aa4e64,64'h317fdb2dface3f77,
64'h1798ff4454da3fa1,64'h10f4d2e8b117c8eb,64'h8b85c27ee4c27a05,64'hfa32e15c4e886138,
64'hb256373e840461ea,64'hfb6921a3de133b8a,64'hed4bdfa524140522,64'h4c740c73ea159d4b,
64'h8ee32067b63a0bb1,64'h70553a9b011648c9,64'h3266a5da6a6edb7d,64'hfffffffefffffff1,
64'h7b13ae612ffa8cba,64'h5a6ea699983d8188,64'hfbd7447e128cbd2f,64'h25fa0114f3b0d464,
64'hff58f19ea0731cd5,64'hcb2345a653affc21,64'h47ea8f0b63c04d38,64'h7bc0e9c9b9f4aafd,
64'h4dba1f70c44a932a,64'h0a3df984fd8d4b60,64'h55281931ab8fc582,64'h65052938d74e90a4,
64'hf58d83521a8cd444,64'h913e1c0a4fafdf66,64'hd84ec4d5cb221841,64'hd212e8cec8a1ed2d,
64'h52bc120e96d36d41,64'hcf1c22e05e886d58,64'hacc3833ef4cf804b,64'h40265167762db5c1,
64'h2ba65b52d7b16755,64'h5e0dbca610ea4244,64'h8613786f669e03bc,64'h5630f7861b6f3d26,
64'h8a571d6878325b67,64'hdcc4194df53c7688,64'hdbe7825afe110978,64'h42cd821357456a45,
64'ha38d268964c594d5,64'hf5aeba1797d9e274,64'h287d4e985b621e77,64'hffffdfff20002001,
64'h31c35693707ff0fd,64'h471db6fa98649a1d,64'h1b5d9404dbf45464,64'h37757208e2a1021b,
64'ha6fa0fe3bfe1caa3,64'h11ba99e61912b7e4,64'h694319b73ad74e57,64'h54ea8dde9bcdf460,
64'hb30249fea3363eb7,64'h10872961a98ab1f8,64'hbb8993978cece8dc,64'h2aa89fc2115650a4,
64'h73885165453beed2,64'h49fceee6592b9b99,64'h96e99e949df66ff4,64'ha4a4eeaf3df82e41,
64'h8907625b5fa6d8f7,64'h4e7f6541087dc789,64'h1fbd6e9f4552731d,64'h8bfed970d671fbb7,
64'hbcc7fa22a6d1fd08,64'h87a6974588be4758,64'h5c2e13fb2613d024,64'hd1970ae9744309b9,
64'h92b1b9f920230f4b,64'hdb490d25f099dc49,64'h6a5efd3020a02909,64'h63a063a150acea56,
64'h77190341b1d05d84,64'h82a9d4db08b24645,64'h93352ed45376dbe7,64'hfffffffeffffff81,
64'hd89d730c7fd465cd,64'hd37534cec1ec0c3e,64'hdeba23f79465e971,64'h2fd008a89d86a31f,
64'hfac78cfc0398e6a1,64'h591a2d389d7fe102,64'h3f54785d1e0269be,64'hde074e50cfa557e5,
64'h6dd0fb882254994e,64'h51efcc27ec6a5b00,64'ha940c98f5c7e2c0e,64'h282949c9ba74851d,
64'hac6c1a97d466a219,64'h89f0e0567d7efb2c,64'hc27626b45910c202,64'h9097467c450f6962,
64'h95e09076b69b6a06,64'h78e11708f4436aba,64'h661c19fca67c0253,64'h01328b3db16dae06,
64'h5d32da97bd8b3aa7,64'hf06de5328752121e,64'h309bc37f34f01ddc,64'hb187bc32db79e92e,
64'h52b8eb47c192db34,64'he620ca75a9e3b43a,64'hdf3c12ddf0884bba,64'h166c109cba2b5226,
64'h1c693450262ca6a3,64'had75d0c3becf1399,64'h43ea74c3db10f3b7,64'hffff000000010001,
64'h8e1ab49c83ff87e7,64'h38edb7d6c324d0e6,64'hdaeca026dfa2a320,64'hbbab9048150810d7,
64'h37d07f22ff0e5513,64'h8dd4cf30c895bf20,64'h4a18cdbcd6ba72b5,64'ha7546ef6de6fa2fe,
64'h98124ffa19b1f5b3,64'h84394b0d4c558fc0,64'hdc4c9cc1676746db,64'h5544fe118ab2851f,
64'h9c428b2d29df768d,64'h4fe77734c95cdcc6,64'hb74cf4a8efb37f9c,64'h2527757eefc17203,
64'h483b12defd36c7b4,64'h73fb2a0a43ee3c46,64'hfdeb74fa2a9398e8,64'h5ff6cb8ab38fddb4,
64'he63fd11a368fe83b,64'h3d34ba3045f23abc,64'he1709fdb309e811e,64'h8cb85751a2184dc2,
64'h958dcfcd01187a54,64'hda48693584cee242,64'h52f7e98405014845,64'h1d031d0d856752ad,
64'hb8c81a108e82ec1d,64'h154ea6dc45923224,64'h99a976a69bb6df34,64'hfffffffefffffc01,
64'hc4eb9869fea32e62,64'h9ba9a67c0f6061ea,64'hf5d11fc2a32f4b82,64'h7e804545ec3518f7,
64'hd63c67e71cc73501,64'hc8d169c6ebff080e,64'hfaa3c2e9f0134def,64'hf03a728c7d2abf22,
64'h6e87dc4412a4ca6d,64'h8f7e61416352d7fe,64'h4a064c7fe3f1606b,64'h414a4e4ed3a428e7,
64'h6360d4c3a33510c3,64'h4f8702b7ebf7d95c,64'h13b135a8c886100a,64'h84ba33e6287b4b0c,
64'haf0483b9b4db502c,64'hc708b84aa21b55cd,64'h30e0cfe833e01295,64'h099459ed8b6d7030,
64'he996d4bfec59d536,64'h836f299b3a9090e9,64'h84de1bfaa780eedf,64'h8c3de19bdbcf496b,
64'h95c75a400c96d99e,64'h310653b44f1da1c9,64'hf9e096f584425dca,64'hb36084e5d15a9130,
64'he349a28131653518,64'h6bae8622f6789cc3,64'h1f53a620d8879db6,64'hfff8000700080001,
64'h70d5a4e81ffc3f34,64'hc76dbeb71926872f,64'hd765013cfd1518fa,64'hdd5c8245a84086b3,
64'hbe83f918f872a897,64'h6ea6798a44adf8fc,64'h50c66de8b5d395a6,64'h3aa377bbf37d17eb,
64'hc0927fd4cd8fad94,64'h21ca586e62ac7dfc,64'he264e6113b3a36d2,64'haa27f08e559428f6,
64'he214596d4efbb464,64'h7f3bb9a84ae6e62e,64'hba67a54c7d9bfcdb,64'h293babf87e0b9017,
64'h41d896f9e9b63d9e,64'h9fd950551f71e22d,64'hef5ba7d8549cc739,64'hffb65c579c7eed9e,
64'h31fe88d8b47f41d1,64'he9a5d1832f91d5df,64'h0b84fee084f408e9,64'h65c2ba9110c26e0c,
64'hac6e7e6c08c3d29c,64'hd24349b22677120a,64'h97bf4c22280a4226,64'he818e86c2b3a9568,
64'hc640d089741760e3,64'haa7536e22c919120,64'hcd4bb538ddb6f99c,64'hfffffffeffffe001,
64'h275cc355f519730a,64'hdd4d33e47b030f4c,64'hae88fe1c197a5c09,64'hf4022a3261a8c7b5,
64'hb1e33f3ee639a802,64'h468b4e3d5ff8406a,64'hd51e1756809a6f71,64'h81d3946ae955f909,
64'h743ee22395265365,64'h7bf30a0f1a96bfec,64'h503264011f8b0356,64'h0a5272789d214736,
64'h1b06a62019a88615,64'h7c3815c15fbecade,64'h9d89ad4644308050,64'h25d19f3543da585c,
64'h78241dd2a6da815b,64'h3845c25b10daae62,64'h87067f429f0094a7,64'h4ca2cf6c5b6b8180,
64'h4cb6a60662cea9a9,64'h1b794cddd4848744,64'h26f0dfd93c0776f4,64'h61ef0ce2de7a4b54,
64'hae3ad20464b6ccec,64'h88329da378ed0e47,64'hcf04b7b32212ee49,64'h9b0427338ad4897b,
64'h1a4d14108b29a8b9,64'h5d74311ab3c4e615,64'hfa9d3106c43cedb0,64'hffc0003f00400001,
64'h86ad2743ffe1f99d,64'h3b6df5bec9343972,64'hbb2809ede8a8c7ca,64'heae4123342043592,
64'hf41fc8ccc39544b3,64'h7533cc55256fc7dd,64'h86336f47ae9cad2e,64'hd51bbde09be8bf57,
64'h0493feac6c7d6c9a,64'h0e52c3741563efdf,64'h13273090d9d1b689,64'h513f8477aca147ab,
64'h10a2cb7177dda319,64'hf9ddcd455737316d,64'hd33d2a68ecdfe6d3,64'h49dd5fc4f05c80b7,
64'h0ec4b7d14db1ecee,64'hfeca82acfb8f1164,64'h7add3ec9a4e639c1,64'hfdb2e2c3e3f76ce9,
64'h8ff446c6a3fa0e87,64'h4d2e8c207c8eaef1,64'h5c27f70427a04748,64'h2e15d48b8613705d,
64'h6373f365461e94db,64'h921a4d9733b8904a,64'hbdfa61154052112c,64'h40c7436859d4ab39,
64'h32068451a0bb0712,64'h53a9b716648c88fb,64'h6a5da9ccedb7ccda,64'hfffffffeffff0001,
64'h3ae61ab0a8cb984f,64'hea699f29d8187a5a,64'h7447f0e5cbd2e043,64'ha011519a0d463da1,
64'h8f19f9fc31cd400b,64'h345a71ecffc2034e,64'ha8f0baba04d37b82,64'h0e9ca35b4aafc844,
64'ha1f7111fa9329b25,64'hdf98507bd4b5ff5d,64'h8193200afc581aae,64'h529393c4e90a39b0,
64'hd8353100cd4430a8,64'he1c0ae0dfdf656ed,64'hec4d6a362184027c,64'h2e8cf9ab1ed2c2df,
64'hc120ee9836d40ad5,64'hc22e12d986d5730f,64'h3833fa18f804a534,64'h65167b64db5c0bfe,
64'h65b5303516754d46,64'hdbca66eea4243a20,64'h3786fecae03bb79f,64'h0f786719f3d25a9d,
64'h71d6902825b6675b,64'h4194ed1fc7687234,64'h7825bd9f10977242,64'hd82139a056a44bd4,
64'hd268a084594d45c8,64'heba188d79e2730a6,64'hd4e9883d21e76d79,64'hfe0001ff02000001,
64'h35693a23ff0fcce4,64'hdb6fadf749a1cb8f,64'hd9404f7445463e4b,64'h572091a11021ac89,
64'ha0fe466d1caa2591,64'ha99e62ac2b7e3ee5,64'h319b7a4174e5696c,64'ha8ddef0adf45fab2,
64'h249ff56363eb64d0,64'h72961ba0ab1f7ef8,64'h99398486ce8db448,64'h89fc23bf650a3d56,
64'h85165b8bbeed18c8,64'hceee6a31b9b98b61,64'h99e9534d66ff3692,64'h4eeafe2982e405b6,
64'h7625be8a6d8f6770,64'hf654156edc788b19,64'hd6e9f6502731ce05,64'hed9716261fbb6741,
64'h7fa236391fd07434,64'h69746105e4757786,64'he13fb8233d023a3e,64'h70aea45d309b82e7,
64'h1b9f9b2d30f4a6d5,64'h90d26cbd9dc4824c,64'hefd308af0290895b,64'h063a1b44cea559c6,
64'h9034228e05d8388f,64'h9d4db8b5246447d6,64'h52ed4e6a6dbe66cd,64'hfffffffefff80001,
64'hd730d586465cc277,64'h534cf955c0c3d2c9,64'ha23f87315e970215,64'h008a8cd56a31ed03,
64'h78cfcfe58e6a0054,64'ha2d38f68fe101a6f,64'h4785d5d5269bdc0b,64'h74e51ada557e4220,
64'h0fb889024994d923,64'hfcc283e4a5affae2,64'h0c99005be2c0d56c,64'h949c9e294851cd7e,
64'hc1a9880c6a21853a,64'h0e057076efb2b761,64'h626b51b80c2013d9,64'h7467cd59f69616f7,
64'h090774c7b6a056a2,64'h117096d236ab9872,64'hc19fd0c8c025299f,64'h28b3db29dae05fed,
64'h2da981abb3aa6a2d,64'hde53377b2121d0fa,64'hbc37f65801ddbcf7,64'h7bc338cf9e92d4e8,
64'h8eb481442db33ad5,64'h0ca769003b43919e,64'hc12decfb84bb920d,64'hc109cd08b5225e9a,
64'h93450428ca6a2e3a,64'h5d0c46c3f1398529,64'ha74c41ef0f3b6bc2,64'hf0000fff10000001,
64'hab49d120f87e671f,64'hdb7d6fc04d0e5c72,64'hca027ba82a31f252,64'hb9048d0a810d6446,
64'h07f2336de5512c83,64'h4cf315665bf1f723,64'h8cdbd20ca72b4b5f,64'h46ef785bfa2fd58b,
64'h24ffab1c1f5b267f,64'h94b0dd0858fbf7bd,64'hc9cc243a746da23c,64'h4fe11dff2851eaac,
64'h28b2dc61f768c63c,64'h77735193cdcc5b02,64'hcf4a9a6f37f9b48c,64'h7757f14e17202dae,
64'hb12df4566c7b3b7d,64'hb2a0ab7de3c458c1,64'hb74fb287398e7022,64'h6cb8b137fddb3a01,
64'hfd11b1cbfe83a19d,64'h4ba3083223abbc2d,64'h09fdc120e811d1e9,64'h857522ec84dc1735,
64'hdcfcd96987a536a8,64'h869365f0ee24125c,64'h7e98457f14844ad1,64'h31d0da26752ace30,
64'h81a114742ec1c474,64'hea6dc5ad23223eac,64'h976a73556df33666,64'hfffffffeffc00001,
64'hb986ac3832e613b2,64'h9a67cab0061e9646,64'h11fc398ff4b810a3,64'h045466ab518f6818,
64'hc67e7f2f7350029d,64'h169c7b4cf080d373,64'h3c2eaeab34dee056,64'ha728d6d5abf210fd,
64'h7dc448124ca6c918,64'he6141f2c2d7fd709,64'h64c802df1606ab60,64'ha4e4f14e428e6bec,
64'h0d4c4069510c29ca,64'h702b83b77d95bb08,64'h135a8dc361009ec5,64'ha33e6ad2b4b0b7b5,
64'h483ba63db502b510,64'h8b84b691b55cc390,64'h0cfe864c01294cf2,64'h459ed94fd702ff67,
64'h6d4c0d5e9d535167,64'hf299bbdf090e87ca,64'he1bfb2c50eede7b3,64'hde19c67ff496a73d,
64'h75a40a256d99d6a4,64'h653b4801da1c8cf0,64'h096f67e225dc9062,64'h084e684ba912f4ca,
64'h9a28214a535171cc,64'he862362189cc2946,64'h3a620f7d79db5e0b,64'h80007fff80000001,
64'h5a4e890cc3f338f3,64'hdbeb7e086872e38a,64'h5013dd47518f928a,64'hc8246859086b222b,
64'h3f919b6f2a896418,64'h6798ab34df8fb916,64'h66de9069395a5af4,64'h377bc2e1d17eac56,
64'h27fd58e1fad933f7,64'ha586e846c7dfbde4,64'h4e6121d9a36d11da,64'h7f08effb428f555e,
64'h4596e310bb4631df,64'hbb9a8ca16e62d80d,64'h7a54d37fbfcda45a,64'hbabf8a73b9016d6d,
64'h896fa2b863d9dbe3,64'h95055bf41e22c603,64'hba7d943ecc73810b,64'h65c589c2eed9d005,
64'he88d8e66f41d0ce1,64'h5d1841931d5de166,64'h4fee0907408e8f48,64'h2ba9176826e0b9a4,
64'he7e6cb523d29b53a,64'h349b2f8b712092dc,64'hf4c22bfba4225685,64'h8e86d134a956717f,
64'h0d08a3a5760e239c,64'h536e2d701911f559,64'hbb539aaf6f99b32c,64'hfffffffefe000001,
64'hcc3561c697309d8b,64'hd33e558430f4b22c,64'h8fe1cc7fa5c08518,64'h22a3355a8c7b40c0,
64'h33f3f9819a8014e2,64'hb4e3da6784069b98,64'he175755aa6f702af,64'h3946b6b25f9087e3,
64'hee224095653648bd,64'h30a0f9686bfeb841,64'h264016fbb0355afd,64'h27278a7714735f5b,
64'h6a62034a88614e50,64'h815c1dbeecadd83d,64'h9ad46e1b0804f628,64'h19f3569aa585bda3,
64'h41dd31efa815a87e,64'h5c25b491aae61c7c,64'h67f43260094a6790,64'h2cf6ca80b817fb36,
64'h6a606af7ea9a8b35,64'h94cddeff48743e49,64'h0dfd962f776f3d91,64'hf0ce3405a4b539e2,
64'had20512e6cceb51d,64'h29da4011d0e4677d,64'h4b7b3f112ee48310,64'h4273425d4897a650,
64'hd1410a569a8b8e5c,64'h4311b1134e614a29,64'hd3107beccedaf057,64'h0004000000000004,
64'hd27448681f99c796,64'hdf5bf04943971c4a,64'h809eea3c8c7c944e,64'h412342ce43591152,
64'hfc8cdb7a544b20bf,64'h3cc559a9fc7dc8ad,64'h36f4834ccad2d79d,64'hbbde170f8bf562af,
64'h3feac710d6c99fb7,64'h2c37423b3efdef1b,64'h73090ecf1b688ece,64'hf8477fdd147aaaed,
64'h2cb71887da318ef6,64'hdcd465107316c063,64'hd2a69c00fe6d22cd,64'hd5fc53a2c80b6b63,
64'h4b7d15c71ecedf14,64'ha82adfa4f1163014,64'hd3eca1fb639c0853,64'h2e2c4e1a76ce8025,
64'h446c733ea0e86701,64'he8c20c9aeaef0b2e,64'h7f70483c04747a3e,64'h5d48bb423705cd1f,
64'h3f365a98e94da9c9,64'ha4d97c5c890496df,64'ha6115fe42112b421,64'h743689a94ab38bf4,
64'h68451d2bb0711ce0,64'h9b716b82c88faac6,64'hda9cd5807ccd995b,64'hfffffffef0000001,
64'h61ab0e3ab984ec52,64'h99f2ac2787a5915a,64'h7f0e64012e0428bc,64'h1519aad563da05ff,
64'h9f9fcc0dd400a70f,64'ha71ed3412034dcbb,64'h0babaadc37b81571,64'hca35b593fc843f17,
64'h711204b229b245e1,64'h8507cb445ff5c207,64'h3200b7de81aad7e7,64'h393c53b9a39afad7,
64'h53101a57430a727d,64'h0ae0edfb656ec1e4,64'hd6a370dc4027b13c,64'hcf9ab4d52c2ded18,
64'h0ee98f7f40ad43ee,64'he12da48f5730e3de,64'h3fa193034a533c7d,64'h67b65406c0bfd9af,
64'h530357c254d459a5,64'ha66ef7fe43a1f244,64'h6fecb17bbb79ec88,64'h8671a03425a9cf09,
64'h690289786675a8e3,64'h4ed2008f87233be7,64'h5bd9f88b7724187e,64'h139a12ec44bd327e,
64'h8a0852bad45c72da,64'h188d889c730a5146,64'h9883df6c76d782b2,64'h0020000000000020,
64'h93a24346fcce3caa,64'hfadf82501cb8e24a,64'h04f751e863e4a26c,64'h091a16741ac88a8e,
64'he466dbd9a25905f1,64'he62acd50e3ee4567,64'hb7a41a675696bce7,64'hdef0b8815fab1573,
64'hff563887b64cfdb7,64'h61ba11daf7ef78d7,64'h9848767bdb44766d,64'hc23bfeefa3d55761,
64'h65b8c43fd18c77af,64'he6a3288998b60312,64'h9534e00df3691662,64'hafe29d1c405b5b12,
64'h5be8ae3af676f89e,64'h4156fd2c88b1809b,64'h9f650fe11ce04292,64'h716270d4b6740127,
64'h236399f707433806,64'h461064de57785969,64'hfb8241e323a3d1ed,64'hea45da13b82e68f6,
64'hf9b2d4c84a6d4e47,64'h26cbe2e94824b6f3,64'h308aff260895a103,64'ha1b44d4d559c5f9d,
64'h4228e9608388e6fd,64'hdb8b5c1a447d562c,64'hd4e6ac09e66ccad2,64'hfffffffe80000001,
64'h0d5871d8cc27628d,64'hcf9561403d2c8acc,64'hf873200c702145dd,64'ha8cd56ab1ed02ff8,
64'hfcfe6072a0053874,64'h38f69a0e01a6e5d3,64'h5d5d56e1bdc0ab88,64'h51adaca5e421f8b2,
64'h889025944d922f05,64'h283e5a26ffae1034,64'h9005bef50d56bf37,64'hc9e29dce1cd7d6b7,
64'h9880d2bc185393e6,64'h57076fdb2b760f20,64'hb51b86e8013d89da,64'h7cd5a6af616f68ba,
64'h774c7bfa056a1f70,64'h096d2481b9871ee9,64'hfd0c981b5299e3e7,64'h3db2a03905fecd75,
64'h981abe14a6a2cd26,64'h3377bff71d0f921b,64'h7f658be0dbcf643d,64'h338d01a52d4e7844,
64'h48144bc633ad4715,64'h7690047e3919df36,64'hdecfc45db920c3ee,64'h9cd0976225e993f0,
64'h504295daa2e396cc,64'hc46c44e398528a30,64'hc41efb67b6bc158c,64'h0100000000000100,
64'h9d121a3be671e54c,64'hd6fc1287e5c71249,64'h27ba8f431f251360,64'h48d0b3a0d6445470,
64'h2336ded412c82f81,64'h31566a8e1f722b31,64'hbd20d33fb4b5e733,64'hf785c410fd58ab92,
64'hfab1c444b267edb1,64'h0dd08edabf7bc6b5,64'hc243b3e2da23b364,64'h11dff7831eaabb02,
64'h2dc622018c63bd75,64'h35194453c5b01889,64'ha9a700739b48b30c,64'h7f14e8e702dad88b,
64'hdf4571d9b3b7c4ee,64'h0ab7e966458c04d6,64'hfb287f0ce702148c,64'h8b1386a8b3a00935,
64'h1b1ccfb93a19c02f,64'h308326f4bbc2cb46,64'hdc120f201d1e8f61,64'h522ed0a4c17347a9,
64'hcd96a649536a7231,64'h365f174b4125b797,64'h8457f93144ad0817,64'h0da26a6face2fce3,
64'h11474b061c4737e6,64'hdc5ae0d823eab15a,64'ha73560553366568a,64'hfffffffb00000001,
64'h6ac38ec6613b1468,64'h7cab0a07e964565a,64'hc399006a810a2ee1,64'h466ab55df6817fbb,
64'he7f3039c0029c399,64'hc7b4d0710d372e97,64'heaeab70fee055c3e,64'h8d6d6531210fc58e,
64'h44812ca66c917824,64'h41f2d138fd70819f,64'h802df7ac6ab5f9b4,64'h4f14ee76e6beb5b2,
64'hc40695e4c29c9f2c,64'hb83b7edb5bb078fe,64'ha8dc374509ec4ecb,64'he6ad357e0b7b45cd,
64'hba63dfd32b50fb7d,64'h4b69240dcc38f748,64'he864c0e194cf1f31,64'hed9501c92ff66ba7,
64'hc0d5f0a93516692c,64'h9bbdffb9e87c90d7,64'hfb2c5f09de7b21e5,64'h9c680d2a6a73c21f,
64'h40a25e339d6a38a6,64'hb48023f4c8cef9ad,64'hf67e22f3c9061f6a,64'he684bb152f4c9f7c,
64'h8214aed7171cb65e,64'h23622722c294517a,64'h20f7db43b5e0ac5a,64'h0800000000000800,
64'he890d1e3338f2a5c,64'hb7e094452e389242,64'h3dd47a19f9289aff,64'h46859d08b222a37e,
64'h19b6f6a196417c07,64'h8ab35471fb915987,64'he9069a02a5af3993,64'hbc2e208eeac55c89,
64'hd58e222c933f6d81,64'h6e8476d5fbde35a8,64'h121d9f1cd11d9b1a,64'h8effbc18f555d810,
64'h6e31100d631deba7,64'ha8ca229f2d80c447,64'h4d3803a1da45985b,64'hf8a7473b16d6c455,
64'hfa2b8ed39dbe276a,64'h55bf4b322c6026b0,64'hd943f86e3810a459,64'h589c35499d0049a4,
64'hd8e67dc9d0ce0178,64'h841937a6de165a2f,64'he0907906e8f47b02,64'h917685280b9a3d46,
64'h6cb532509b539182,64'hb2f8ba5b092dbcb7,64'h22bfc98e256840b4,64'h6d13537d6717e718,
64'h8a3a5830e239bf30,64'he2d706c71f558aca,64'h39ab02ae9b32b44b,64'hffffffdf00000001,
64'h561c763609d8a33d,64'he55850424b22b2cd,64'h1cc8035a08517702,64'h3355aaf1b40bfdd6,
64'h3f981ce7014e1cc1,64'h3da6838e69b974b2,64'h5755b886702ae1e9,64'h6b6b298d087e2c6c,
64'h24096535648bc11e,64'h0f9689c9eb840cf6,64'h016fbd6755afcd9c,64'h78a773b935f5ad8e,
64'h2034af2c14e4f95a,64'hc1dbf6dfdd83c7eb,64'h46e1ba2d4f627653,64'h3569abf75bda2e61,
64'hd31efe9e5a87dbe3,64'h5b49207061c7ba3e,64'h43260713a678f981,64'h6ca80e507fb35d31,
64'h06af854fa8b3495a,64'hddeffdd343e486b4,64'hd962f855f3d90f21,64'he3406957539e10f4,
64'h0512f19eeb51c52e,64'ha4011fab4677cd63,64'hb3f117a54830fb49,64'h3425d8b07a64fbd9,
64'h10a576bcb8e5b2ec,64'h1b11391714a28bcf,64'h07beda1eaf0562cf,64'h4000000000004000,
64'h44868f209c7952d9,64'hbf04a22e71c4920b,64'heea3d0d0c944d7f7,64'h342ce84791151bee,
64'hcdb7b50cb20be038,64'h559aa393dc8acc34,64'h4834d01c2d79cc91,64'he171047c562ae443,
64'hac71116a99fb6c02,64'h7423b6b2def1ad3d,64'h90ecf8e688ecd8d0,64'h77fde0cbaaaec07c,
64'h7188806e18ef5d35,64'h465114fe6c062233,64'h69c01d10d22cc2d6,64'hc53a39dfb6b622a1,
64'hd15c76a3edf13b49,64'hadfa59936301357e,64'hca1fc377c08522c2,64'hc4e1aa4ee8024d1e,
64'hc733ee5486700bba,64'h20c9bd3af0b2d174,64'h0483c83e47a3d809,64'h8bb429445cd1ea2c,
64'h65a99287da9c8c0d,64'h97c5d2dd496de5b3,64'h15fe4c722b42059f,64'h689a9bee38bf38bd,
64'h51d2c18b11cdf97c,64'h16b8363ffaac5649,64'hcd581575d995a257,64'hfffffeff00000001,
64'hb0e3b1b24ec519e6,64'h2ac2821959159661,64'he6401ad0428bb810,64'h9aad578ea05feeaf,
64'hfcc0e7390a70e607,64'hed341c744dcba58f,64'hbaadc43581570f46,64'h5b594c6b43f1635d,
64'h204b29ac245e08ef,64'h7cb44e4f5c2067b0,64'h0b7deb3aad7e6ce0,64'hc53b9dccafad6c6d,
64'h01a57961a727cacf,64'h0edfb704ec1e3f52,64'h370dd16c7b13b296,64'hab4d5fbbded17307,
64'h98f7f4f8d43edf12,64'hda4903850e3dd1ee,64'h1930389f33c7cc06,64'h65407286fd9ae985,
64'h357c2a7d459a4ad0,64'hef7feea01f24359a,64'hcb17c2b59ec87902,64'h1a034ac19cf08799,
64'h28978cf75a8e2970,64'h2008fd5f33be6b13,64'h9f88bd2f4187da43,64'ha12ec584d327dec7,
64'h852bb5e5c72d9760,64'hd889c8b8a5145e78,64'h3df6d0f5782b1678,64'h000000020001fffe,
64'h24347906e3ca96c6,64'hf82511788e249053,64'h751e868d4a26bfb1,64'ha167423d88a8df6f,
64'h6dbda86b905f01ba,64'hacd51ca0e456619e,64'h41a680e36bce6486,64'h0b8823e9b1572211,
64'h63888b59cfdb600b,64'ha11db599f78d69e5,64'h8767c7384766c67c,64'hbfef0660557603dd,
64'h8c440373c77ae9a5,64'h3288a7f560311196,64'h4e00e889916616ad,64'h29d1cf03b5b11502,
64'h8ae3b5256f89da42,64'h6fd2cca01809abeb,64'h50fe1bc40429160a,64'h270d527d401268ea,
64'h399f72aa33805dca,64'h064de9d885968b9f,64'h241e41f23d1ec048,64'h5da14a26e68f515c,
64'h2d4c9441d4e46065,64'hbe2e96ee4b6f2d94,64'haff263915a102cf8,64'h44d4df74c5f9c5e5,
64'h8e960c5a8e6fcbde,64'hb5c1b1ffd562b248,64'h6ac0abb4ccad12b2,64'hfffff7ff00000001,
64'h871d8d977628cf2b,64'h561410cbc8acb307,64'h3200d689145dc079,64'hd56abc7902ff7574,
64'he60739cf53873031,64'h69a0e3a96e5d2c71,64'hd56e21b10ab87a2b,64'hdaca635c1f8b1ae6,
64'h02594d6222f04777,64'he5a2727de1033d7d,64'h5bef59d56bf36700,64'h29dcee6b7d6b6362,
64'h0d2bcb0d393e5678,64'h76fdb82760f1fa90,64'hb86e8b64d89d94af,64'h5a6afde3f68b9833,
64'hc7bfa7caa1f6f88c,64'hd2481c2e71ee8f6a,64'hc981c4f99e3e6030,64'h2a03943aecd74c25,
64'habe153eb2cd2567f,64'h7bff7507f921acc9,64'h58be15b2f643c80a,64'hd01a560ce7843cc8,
64'h44bc67bbd4714b7f,64'h0047eafa9df35897,64'hfc45e97e0c3ed214,64'h09762c2b993ef633,
64'h295daf32396cbafc,64'hc44e45cb28a2f3ba,64'hefb687acc158b3bf,64'h00000010000ffff0,
64'h21a3c8381e54b62f,64'hc1288bcb71248291,64'ha8f4346d5135fd85,64'h0b3a11f14546fb73,
64'h6ded435f82f80dcd,64'h66a8e50c22b30ceb,64'h0d34071d5e73242e,64'h5c411f4d8ab91088,
64'h1c445ad17edb0055,64'h08edacd4bc6b4f23,64'h3b3e39c63b3633dc,64'hff783307abb01ee3,
64'h62201ba23bd74d24,64'h94453fac01888caf,64'h7007444e8b30b566,64'h4e8e781ead88a80f,
64'h571da92f7c4ed20c,64'h7e966503c04d5f55,64'h87f0de222148b04e,64'h386a93eb0093474f,
64'hccfb95529c02ee4f,64'h326f4ec42cb45cf8,64'h20f20f92e8f6023f,64'hed0a5139347a8ade,
64'h6a64a20fa7230327,64'hf174b7775b796c9b,64'h7f931c8fd08167bb,64'h26a6fba82fce2f26,
64'h74b062d8737e5eec,64'hae0d9003ab15923b,64'h56055da96568958d,64'hffffbfff00000001,
64'h38ec6cbfb1467954,64'hb0a0866045659836,64'h9006b449a2ee03c7,64'hab55e3ce17fbab9a,
64'h3039ce819c398181,64'h4d071d4e72e96385,64'hab710d8e55c3d152,64'hd6531ae6fc58d72a,
64'h12ca6b1117823bb8,64'h2d1393f60819ebe1,64'hdf7acead5f9b37fe,64'h4ee7735ceb5b1b0f,
64'h695e5869c9f2b3c0,64'hb7edc13e078fd47d,64'hc3745b2bc4eca573,64'hd357ef21b45cc196,
64'h3dfd3e5b0fb7c45a,64'h9240e1798f747b4a,64'h4c0e27d2f1f3017a,64'h501ca1d866ba6127,
64'h5f0a9f5e6692b3f3,64'hdffba842c90d6645,64'hc5f0ad99b21e404e,64'h80d2b06d3c21e63a,
64'h25e33de0a38a5bf6,64'h023f57d4ef9ac4b8,64'he22f4bf761f69099,64'h4bb1615cc9f7b198,
64'h4aed7992cb65d7df,64'h22722e5f45179dca,64'h7db43d6d0ac59df1,64'h00000080007fff80,
64'h0d1e41c1f2a5b177,64'h09445e6189241482,64'h47a1a36f89afec23,64'h59d08f8a2a37db98,
64'h6f6a1aff17c06e65,64'h3547286415986755,64'h69a038eaf3992170,64'he208fa6e55c8843e,
64'he222d68bf6d802a8,64'h476d66a5e35a7918,64'hd9f1ce32d9b19edf,64'hfbc198445d80f711,
64'h1100dd14deba691d,64'ha229fd640c446574,64'h803a22775985ab2d,64'h7473c0f76c454076,
64'hb8ed497de276905e,64'hf4b32821026afaa5,64'h3f86f1150a45826c,64'hc3549f59049a3a77,
64'h67dcaa9ae0177272,64'h937a762265a2e7bf,64'h07907c9847b011f7,64'h685289d0a3d456e9,
64'h5325108039181935,64'h8ba5bbc1dbcb64d1,64'hfc98e481840b3dd5,64'h3537dd427e71792f,
64'ha58316c69bf2f75d,64'h706c802258ac91d3,64'hb02aed4d2b44ac66,64'hfffdffff00000001,
64'hc76365fe8a33ca9f,64'h850433072b2cc1ab,64'h8035a25117701e34,64'h5aaf1e75bfdd5ccb,
64'h81ce740de1cc0c07,64'h6838ea75974b1c26,64'h5b886c77ae1e8a8b,64'hb298d73de2c6b94a,
64'h96535888bc11ddc0,64'h689c9fb140cf5f07,64'hfbd67570fcd9bfea,64'h773b9ae95ad8d876,
64'h4af2c3514f959dfd,64'hbf6e09f53c7ea3e3,64'h1ba2d96427652b92,64'h9abf7913a2e60caa,
64'hefe9f2d97dbe22cf,64'h92070bd07ba3da4c,64'h60713e998f980bce,64'h80e50ec535d30936,
64'hf854faf534959f96,64'hffdd421c486b3222,64'h2f856cd390f2026a,64'h0695836de10f31cc,
64'h2f19ef061c52dfaf,64'h11fabea77cd625c0,64'h117a5fc20fb484c1,64'h5d8b0ae84fbd8cbe,
64'h576bcc985b2ebef6,64'h139172fb28bcee4f,64'heda1eb6b562cef85,64'h0000040003fffc00,
64'h68f20e0f952d8bb8,64'h4a22f30c4920a410,64'h3d0d1b7e4d7f6116,64'hce847c5351bedcbe,
64'h7b50d7fbbe037325,64'haa394321acc33aa7,64'h4d01c75a9cc90b7d,64'h1047d379ae4421e9,
64'h1116b466b6c01539,64'h3b6b35311ad3c8be,64'hcf8e719ccd8cf6f2,64'hde0cc229ec07b881,
64'h8806e8a6f5d348e8,64'h114feb2562232b9b,64'h01d113becc2d5964,64'ha39e07be622a03ad,
64'hc76a4bf413b482eb,64'ha599410f1357d521,64'hfc3788a9522c135f,64'h1aa4face24d1d3b2,
64'h3ee554da00bb938d,64'h9bd3b1172d173df4,64'h3c83e4c23d808fb8,64'h42944e881ea2b745,
64'h99288403c8c0c9a6,64'h5d2dde12de5b2684,64'he4c724132059eea1,64'ha9beea14f38bc977,
64'h2c18b639df97bae3,64'h83640115c5648e95,64'h81576a6e5a25632b,64'hffefffff00000001,
64'h3b1b2ffa519e54f2,64'h2821983d59660d54,64'h01ad128cbb80f19c,64'hd578f3affeeae656,
64'h0e73a0730e606034,64'h41c753afba58e12d,64'hdc4363bf70f45456,64'h94c6b9f41635ca4b,
64'hb29ac449e08eedfc,64'h44e4fd8d067af835,64'hdeb3ab8ee6cdff49,64'hb9dcd74dd6c6c3ad,
64'h57961a8c7cacefe6,64'hfb704faee3f51f13,64'hdd16cb213b295c90,64'hd5fbc8a11730654c,
64'h7f4f96d2edf11671,64'h90385e87dd1ed25c,64'h0389f4cf7cc05e6d,64'h0728762dae9849ac,
64'hc2a7d7b0a4acfca9,64'hfeea10e943599109,64'h7c2b669d8790134f,64'h34ac1b6f08798e60,
64'h78cf7831e296fd77,64'h8fd5f53be6b12e00,64'h8bd2fe107da42608,64'hec5857447dec65ee,
64'hbb5e64c4d975f7ae,64'h9c8b97d945e77278,64'h6d0f5b61b1677c21,64'h000020001fffe000,
64'h4790707fa96c5dbd,64'h511798644905207e,64'he868dbf36bfb08af,64'h7423e2a08df6e5ea,
64'hda86bfe0f01b9925,64'h51ca19126619d533,64'h680e3ad6e6485be6,64'h823e9bcd72210f48,
64'h88b5a335b600a9c8,64'hdb59a989d69e45ef,64'h7c738cec6c67b78a,64'hf0661155603dc402,
64'h4037453bae9a473c,64'h8a7f592b11195cd8,64'h0e889df6616acb20,64'h1cf03df811501d63,
64'h3b525fa69da41752,64'h2cca087d9abea903,64'he1bc455191609af1,64'hd527d671268e9d90,
64'hf72aa6d105dc9c67,64'hde9d88bd68b9ef9c,64'he41f2612ec047dbf,64'h14a27442f515ba26,
64'hc944202246064d2c,64'he96ef098f2d9341e,64'h263920a002cf7501,64'h4df750ac9c5e4bb3,
64'h60c5b1cffcbdd717,64'h1b2008b22b2474a4,64'h0abb5376d12b1954,64'hff7fffff00000001,
64'hd8d97fd38cf2a78f,64'h410cc1ebcb306a9f,64'h0d689465dc078ce0,64'habc79d85f75732aa,
64'h739d0398730301a0,64'h0e3a9d7fd2c70966,64'he21b1e0187a2a2aa,64'ha635cfa4b1ae5254,
64'h94d6225404776fdb,64'h2727ec6a33d7c1a6,64'hf59d5c7d366ffa42,64'hcee6ba73b6361d63,
64'hbcb0d465e5677f2e,64'hdb827d7e1fa8f891,64'he8b6590fd94ae47a,64'hafde450eb9832a5a,
64'hfa7cb69a6f88b385,64'h81c2f442e8f692dc,64'h1c4fa67be602f368,64'h3943b16d74c24d60,
64'h153ebd8b2567e542,64'hf75087511acc8841,64'he15b34ef3c809a75,64'ha560db7943cc72ff,
64'hc67bc19214b7ebb5,64'h7eafa9e335896ffc,64'h5e97f087ed21303c,64'h62c2ba2aef632f69,
64'hdaf3262bcbafbd6b,64'he45cbece2f3b93bc,64'h687adb108b3be105,64'h00010000ffff0000,
64'h3c8383ff4b62ede6,64'h88bcc324482903ee,64'h4346dfa25fd84571,64'ha11f15076fb72f4d,
64'hd435ff0d80dcc922,64'h8e50c89530cea996,64'h4071d6ba3242df2d,64'h11f4de6f91087a3c,
64'h45ad19b1b0054e3c,64'hdacd4c54b4f22f72,64'he39c6766633dbc4d,64'h83308ab201ee2009,
64'h01ba29df74d239de,64'h53fac95c88cae6bc,64'h7444efb30b565900,64'he781efc08a80eb18,
64'hda92fd35ed20ba8f,64'h665043edd5f54817,64'h0de22a938b04d781,64'ha93eb38f3474ec7a,
64'hb955368f2ee4e331,64'hf4ec45f145cf7cda,64'h20f9309e6023edf1,64'ha513a217a8add130,
64'h4a2101183032695a,64'h4b7784ce96c9a0e9,64'h31c90501167ba807,64'h6fba8566e2f25d96,
64'h062d8e82e5eeb8b5,64'hd90045915923a520,64'h55da9bb68958caa0,64'hfbffffff00000001,
64'hc6cbfea267953c72,64'h08660f60598354f6,64'h6b44a32ee03c6700,64'h5e3cec34bab9954b,
64'h9ce81cc698180cfd,64'h71d4ebfe96384b30,64'h10d8f0133d151549,64'h31ae7d2a8d72929b,
64'ha6b112a423bb7ed4,64'h393f63529ebe0d2f,64'haceae3f0b37fd209,64'h7735d3a3b1b0eb12,
64'he586a3342b3bf96b,64'hdc13ebf6fd47c482,64'h45b2c885ca5723c9,64'h7ef2287acc1952cb,
64'hd3e5b4da7c459c21,64'h0e17a21b47b496dc,64'he27d33df30179b40,64'hca1d8b6ca6126aff,
64'ha9f5ec592b3f2a10,64'hba843a8fd6644201,64'h0ad9a780e404d3a1,64'h2b06dbcf1e6397f3,
64'h33de0c96a5bf5da2,64'hf57d4f1cac4b7fdd,64'hf4bf8441690981de,64'h1615d15a7b197b45,
64'hd79931645d7deb52,64'h22e5f67879dc9dd9,64'h43d6d88759df0825,64'h00080007fff80000,
64'he41c1ffb5b176f2f,64'h45e6192641481f6c,64'h1a36fd14fec22b86,64'h08f8a8407db97a63,
64'ha1aff87206e6490a,64'h728644ad86754cac,64'h038eb5d39216f966,64'h8fa6f37c8843d1e0,
64'h2d68cd8f802a71de,64'hd66a62aba7917b8a,64'h1ce33b3a19ede261,64'h198455940f710044,
64'h0dd14efba691cef0,64'h9fd64ae6465735de,64'ha2277d9b5ab2c7fd,64'h3c0f7e0b540758b9,
64'hd497e9b56905d472,64'h32821f71afaa40b5,64'h6f11549c5826bc08,64'h49f59c7ea3a763cb,
64'hcaa9b47e77271983,64'ha7622f912e7be6c9,64'h07c984f4011f6f87,64'h289d10c2456e897b,
64'h510808c381934ace,64'h5bbc2676b64d0746,64'h8e482809b3dd4037,64'h7dd42b3a1792ecad,
64'h316c74172f75c5a8,64'hc8022c90c91d28fa,64'haed4ddb64ac654fe,64'hdfffffff00000001,
64'h365ff5193ca9e38a,64'h43307b02cc1aa7b0,64'h5a25197a01e337fd,64'hf1e761a7d5ccaa56,
64'he740e638c0c067e4,64'h8ea75ff7b1c2597d,64'h86c78099e8a8aa48,64'h8d73e9556b9494d7,
64'h358895261ddbf69b,64'hc9fb1a95f5f06977,64'h67571f8a9bfe9043,64'hb9ae9d208d87588d,
64'h2c3519a859dfcb51,64'he09f5fbdea3e240a,64'h2d96443052b91e46,64'hf79143d960ca9655,
64'h9f2da6d9e22ce102,64'h70bd10da3da4b6e0,64'h13e99f0080bcd9f9,64'h50ec5b6b309357f2,
64'h4faf62ce59f9507b,64'hd421d483b3221003,64'h56cd3c0720269d08,64'h5836de79f31cbf97,
64'h9ef064b62dfaed0f,64'habea78ec625bfee1,64'ha5fc2212484c0ee9,64'hb0ae8ad3d8cbda28,
64'hbcc98b28ebef5a8a,64'h172fb3c4cee4eec7,64'h1eb6c43ccef84126,64'h0040003fffc00000,
64'h20e0ffe1d8bb7971,64'h2f30c9340a40fb5e,64'hd1b7e8a7f6115c30,64'h47c54203edcbd318,
64'h0d7fc3953732484b,64'h9432256f33aa655d,64'h1c75ae9c90b7cb30,64'h7d379be8421e8efc,
64'h6b466c7d01538eef,64'hb35315633c8bdc4a,64'he719d9d0cf6f1308,64'hcc22aca07b880220,
64'h6e8a77dd348e7780,64'hfeb2573632b9aeec,64'h113becdfd5963fe3,64'he07bf05ba03ac5c7,
64'ha4bf4db1482ea38a,64'h9410fb8e7d5205a7,64'h788aa4e5c135e03d,64'h4face3f71d3b1e56,
64'h554da3f9b938cc12,64'h3b117c8e73df3643,64'h3e4c27a008fb7c38,64'h44e886132b744bd7,
64'h8840461e0c9a566e,64'hdde133b7b2683a2e,64'h724140519eea01b4,64'heea159d3bc976565,
64'h8b63a0ba7bae2d3f,64'h4011648c48e947ca,64'h76a6edb75632a7eb,64'hfffffffe00000002,
64'hb2ffa8cae54f1c4f,64'h1983d81860d53d7e,64'hd128cbd20f19bfe6,64'h8f3b0d45ae6552a9,
64'h3a0731cd06033f19,64'h753affc18e12cbe4,64'h363c04d34545523c,64'h6b9f4aaf5ca4a6b4,
64'hac44a931eedfb4d7,64'h4fd8d4b5af834bb2,64'h3ab8fc57dff48215,64'hcd74e9096c3ac463,
64'h61a8cd43cefe5a87,64'h04fafdf651f12049,64'h6cb2218395c8f22f,64'hbc8a1ed20654b2a1,
64'hf96d36d31167080c,64'h85e886d4ed25b6fd,64'h9f4cf80405e6cfc8,64'h8762db5b849abf8e,
64'h7d7b1674cfca83d6,64'ha10ea42399108012,64'hb669e03b0134e83e,64'hc1b6f3d198e5fcb6,
64'hf78325b56fd76874,64'h5f53c76812dff703,64'h2fe1109742607743,64'h857456a3c65ed13b,
64'he64c594c5f7ad44b,64'hb97d9e2677277638,64'hf5b621e677c20930,64'h020001fffe000000,
64'h0707ff0fc5dbcb87,64'h798649a15207daef,64'h8dbf4545b08ae17a,64'h3e2a10216e5e98be,
64'h6bfe1ca9b9924258,64'ha1912b7d9d532ae4,64'he3ad74e485be5980,64'he9bcdf4510f477dd,
64'h5a3363eb0a9c7775,64'h9a98ab1ee45ee24b,64'h38cece8d7b789839,64'h61156509dc4010fa,
64'h7453beeca473bbfd,64'hf592b9b895cd7759,64'h89df66feacb1ff18,64'h03df82e401d62e31,
64'h25fa6d8f41751c4b,64'ha087dc77ea902d34,64'hc455273109af01e5,64'h7d671fbae9d8f2ae,
64'haa6d1fcfc9c6608e,64'hd88be4749ef9b217,64'hf2613d0147dbe1bf,64'h2744309b5ba25eb6,
64'h420230f464d2b36c,64'hef099dc39341d16a,64'h920a028ff7500d9d,64'h750acea4e4bb2b21,
64'h5b1d05d7dd7169f4,64'h008b2464474a3e4e,64'hb5376dbdb1953f55,64'hfffffff700000009,
64'h97fd465c2a78e273,64'hcc1ec0c306a9ebf0,64'h89465e9678cdff2a,64'h79d86a31732a9544,
64'hd0398e693019f8c7,64'ha9d7fe0f70965f1d,64'hb1e0269b2a2a91df,64'h5cfa557de525359d,
64'h6225499476fda6b3,64'h7ec6a5af7c1a5d8e,64'hd5c7e2bfffa410a7,64'h6ba7485161d62312,
64'h0d466a2177f2d435,64'h27d7efb28f890248,64'h65910c1fae479175,64'he450f69532a59503,
64'hcb69b69f8b384059,64'h2f4436ab692db7e4,64'hfa67c0242f367e3c,64'h3b16dae024d5fc6c,
64'hebd8b3a97e541ead,64'h08752121c884008b,64'hb34f01dd09a741eb,64'h0db79e92c72fe5aa,
64'hbc192db27ebb4399,64'hfa9e3b4296ffb816,64'h7f0884bb1303ba17,64'h2ba2b52232f689d4,
64'h3262ca69fbd6a251,64'hcbecf138b93bb1bb,64'hadb10f3abe104979,64'h10000ffff0000000,
64'h383ff87e2ede5c38,64'hcc324d0d903ed775,64'h6dfa2a3184570bcc,64'hf150810c72f4c5ef,
64'h5ff0e550cc9212bd,64'h0c895bf1ea99571b,64'h1d6ba72b2df2cbf9,64'h4de6fa2f87a3bee1,
64'hd19b1f5a54e3bba6,64'hd4c558fb22f71254,64'hc676746cdbc4c1c7,64'h08ab2851e20087cd,
64'ha29df768239ddfe5,64'hac95cdcbae6bbac1,64'h4efb37f9658ff8bc,64'h1efc17200eb17188,
64'h2fd36c7b0ba8e257,64'h043ee3c45481699b,64'h22a9398e4d780f22,64'heb38fdda4ec7956d,
64'h5368fe834e33046b,64'hc45f23aaf7cd90b2,64'h9309e8113edf0df1,64'h3a2184dbdd12f5af,
64'h101187a526959b5e,64'h784cee239a0e8b49,64'h90501483ba806ce4,64'ha856752a25d95905,
64'hd8e82ec0eb8b4f9e,64'h045923223a51f270,64'ha9bb6df28ca9faa3,64'hffffffbf00000041,
64'hbfea32e553c71394,64'h60f6061e354f5f7a,64'h4a32f4b7c66ff94c,64'hcec3518e9954aa1d,
64'h81cc734f80cfc632,64'h4ebff08084b2f8e3,64'h8f0134de51548ef3,64'he7d2abf12929ace6,
64'h112a4ca6b7ed3595,64'hf6352d7ee0d2ec6d,64'hae3f1605fd208532,64'h5d3a428e0eb1188d,
64'h6a33510bbf96a1a8,64'h3ebf7d957c48123f,64'h2c886100723c8ba5,64'h2287b4b0952ca811,
64'h5b4db50259c202c2,64'h7a21b55c496dbf1f,64'hd33e012879b3f1d9,64'hd8b6d70226afe35f,
64'h5ec59d52f2a0f561,64'h43a9090e44200458,64'h9a780eed4d3a0f53,64'h6dbcf496397f2d50,
64'he0c96d98f5da1cc3,64'hd4f1da1bb7fdc0a9,64'hf84425db981dd0b5,64'h5d15a91297b44e9f,
64'h93165350deb51287,64'h5f6789cbc9dd8dd2,64'h6d8879daf0824bc3,64'h80007fff80000000,
64'hc1ffc3f276f2e1bf,64'h6192687281f6bba2,64'h6fd1518f22b85e5d,64'h8a84086a97a62f71,
64'hff872a88649095e6,64'h644adf8f54cab8d8,64'heb5d39596f965fc8,64'h6f37d17e3d1df706,
64'h8cd8fad8a71ddd2a,64'ha62ac7df17b8929a,64'h33b3a36cde260e32,64'h4559428f10043e68,
64'h14efbb461ceeff23,64'h64ae6e62735dd603,64'h77d9bfcd2c7fc5de,64'hf7e0b900758b8c40,
64'h7e9b63d95d4712b7,64'h21f71e22a40b4cd8,64'h1549cc736bc0790f,64'h59c7eed9763cab61,
64'h9b47f41c71982356,64'h22f91d5dbe6c858a,64'h984f408df6f86f84,64'hd10c26dfe897ad77,
64'h808c3d2934acdaf0,64'hc267711fd0745a45,64'h8280a421d403671c,64'h42b3a9562ecac823,
64'hc741760d5c5a7cea,64'h22c91911d28f9380,64'h4ddb6f99654fd513,64'hfffffdff00000201,
64'hff51972f9e389c9b,64'h07b030f4aa7afbcd,64'h5197a5c0337fca5e,64'h761a8c7acaa550e2,
64'h0e639a80067e318c,64'h75ff84062597c716,64'h7809a6f68aa47794,64'h3e955f90494d6729,
64'h89526535bf69aca8,64'hb1a96bfe06976361,64'h71f8b034e904298b,64'he9d214727588c466,
64'h519a8860fcb50d3d,64'hf5fbecace24091f7,64'h6443080491e45d27,64'h143da585a9654087,
64'hda6da814ce10160e,64'hd10daae54b6df8f5,64'h99f00949cd9f8ec2,64'hc5b6b817357f1af2,
64'hf62cea999507ab06,64'h1d484874210022be,64'hd3c0776e69d07a94,64'h6de7a4b4cbf96a7d,
64'h064b6cceaed0e611,64'ha78ed0e3bfee0542,64'hc2212ee3c0ee85a1,64'he8ad4896bda274f6,
64'h98b29a8af5a89434,64'hfb3c4e604eec6e8e,64'h6c43ceda84125e15,64'h0003fffffffffffc,
64'h0ffe1f99b7970df2,64'h0c9343970fb5dd0d,64'h7e8a8c7c15c2f2e5,64'h54204358bd317b84,
64'hfc39544a2484af29,64'h2256fc7da655c6bd,64'h5ae9cad27cb2fe39,64'h79be8bf4e8efb82d,
64'h66c7d6c938eee94c,64'h31563efdbdc494cb,64'h9d9d1b67f130718f,64'h2aca147a8021f33e,
64'ha77dda30e777f918,64'h257373169aeeb015,64'hbecdfe6c63fe2eed,64'hbf05c80aac5c61f9,
64'hf4db1ecdea3895b5,64'h0fb8f116205a66bf,64'haa4e639b5e03c878,64'hce3f76cdb1e55b06,
64'hda3fa0e78cc11aac,64'h17c8eaeef3642c4f,64'hc27a0473b7c37c1c,64'h8861370544bd6bb2,
64'h0461e94da566d77c,64'h133b890483a2d222,64'h14052112a01b38dc,64'h159d4ab376564116,
64'h3a0bb070e2d3e74a,64'h1648c88f947c9bff,64'h6edb7ccd2a7ea896,64'hffffefff00001001,
64'hfa8cb983f1c4e4d1,64'h3d8187a553d7de68,64'h8cbd2e039bfe52ee,64'hb0d463d9552a870d,
64'h731cd40033f18c60,64'haffc20342cbe38ad,64'hc04d37b75523bc9d,64'hf4aafc834a6b3947,
64'h4a9329b1fb4d653c,64'h8d4b5ff534bb1b03,64'h8fc581aa48214c55,64'h4e90a39aac462329,
64'h8cd44309e5a869e6,64'hafdf656e12048fb1,64'h221840278f22e935,64'ha1ed2c2d4b2a0438,
64'hd36d40ac7080b06a,64'h886d57305b6fc7a2,64'hcf804a526cfc760c,64'h2db5c0bfabf8d78a,
64'hb16754d3a83d5829,64'hea4243a1080115f0,64'h9e03bb794e83d49a,64'h6f3d25a95fcb53e5,
64'h325b667576873088,64'h3c768722ff702a0b,64'h1109772407742d02,64'h456a44bced13a7a9,
64'hc594d45bad44a19c,64'hd9e2730977637469,64'h621e76d72092f0a5,64'h001fffffffffffe0,
64'h7ff0fccdbcb86f90,64'h649a1cb87daee868,64'hf45463e3ae179725,64'ha1021ac7e98bdc1e,
64'he1caa25824257941,64'h12b7e3ee32ae35e7,64'hd74e5695e597f1c6,64'hcdf45faa477dc165,
64'h363eb64cc7774a5d,64'h8ab1f7eeee24a657,64'hece8db4389838c74,64'h5650a3d5010f99ef,
64'h3beed18c3bbfc8bb,64'h2b9b98b5d77580a7,64'hf66ff3681ff17763,64'hf82e405a62e30fc3,
64'ha6d8f67651c4ada1,64'h7dc788b102d335f8,64'h52731cdff01e43bb,64'h71fbb6738f2ad82a,
64'hd1fd07426608d55a,64'hbe4757779b216278,64'h13d023a3be1be0da,64'h4309b82e25eb5d8c,
64'h230f4a6d2b36bbe0,64'h99dc48241d169110,64'ha029089500d9c6e0,64'hacea559bb2b208b0,
64'hd05d8388169f3a4f,64'hb246447ca3e4dff8,64'h76dbe66c53f544ad,64'hffff7fff00008001,
64'hd465cc268e272681,64'hec0c3d2b9ebef33f,64'h65e97020dff2976c,64'h86a31ecfa9543863,
64'h98e6a0049f8c62fd,64'h7fe101a665f1c563,64'h0269bdc0a91de4e2,64'ha557e4215359ca31,
64'h54994d91da6b29de,64'h6a5affada5d8d814,64'h7e2c0d56410a62a4,64'h74851cd762311946,
64'h66a218532d434f2c,64'h7efb2b7590247d83,64'h10c2013d791749a7,64'h0f69616f595021bb,
64'h9b6a05698405834a,64'h436ab986db7e3d0c,64'h7c02529967e3b05a,64'h6dae05fe5fc6bc4f,
64'h8b3aa6a241eac143,64'h52121d0f4008af79,64'hf01ddbce741ea4cc,64'h79e92d4dfe5a9f25,
64'h92db33acb439843f,64'he3b43918fb815057,64'h884bb9203ba16810,64'h2b5225e9689d3d46,
64'h2ca6a2e36a250cda,64'hcf139851bb1ba342,64'h10f3b6bc04978525,64'h00ffffffffffff00,
64'hff87e670e5c37c7d,64'h24d0e5c6ed77433d,64'ha2a31f2470bcb921,64'h0810d6444c5ee0eb,
64'h0e5512c8212bca01,64'h95bf1f719571af38,64'hba72b4b52cbf8e2a,64'h6fa2fd583bee0b22,
64'hb1f5b2673bba52e7,64'h558fbf7b712532b4,64'h6746da234c1c6399,64'hb2851eaa087ccf76,
64'hdf768c62ddfe45d7,64'h5cdcc5afbbac0537,64'hb37f9b47ff8bbb11,64'hc17202da17187e11,
64'h36c7b3b78e256d03,64'hee3c458b1699afbd,64'h9398e70180f21dd6,64'h8fddb39f7956c14d,
64'h8fe83a193046aaca,64'hf23abbc1d90b13bb,64'h9e811d1df0df06d0,64'h184dc1732f5aec5e,
64'h187a536a59b5deff,64'hcee24124e8b4887c,64'h014844ad06ce36fb,64'h6752ace29590457b,
64'h82ec1c46b4f9d272,64'h923223ea1f26ffbb,64'hb6df33659faa2565,64'hfffbffff00040001,
64'ha32e613a71393402,64'h6061e963f5f799f1,64'h2f4b8109ff94bb5d,64'h3518f6814aa1c314,
64'hc7350028fc6317e4,64'hff080d362f8e2b15,64'h134dee0548ef2710,64'h2abf210f9ace5183,
64'ha4ca6c90d3594eee,64'h52d7fd702ec6c09d,64'hf1606ab50853151d,64'ha428e6be1188ca2d,
64'h3510c29c6a1a795d,64'hf7d95baf8123ec15,64'h861009ebc8ba4d38,64'h7b4b0b7aca810dd8,
64'hdb502b50202c1a4c,64'h1b55cc38dbf1e85e,64'he01294ce3f1d82cd,64'h6d702ff5fe35e275,
64'h59d535160f560a14,64'h9090e87c00457bc6,64'h80eede7aa0f52659,64'hcf496a72f2d4f925,
64'h96d99d69a1cc21f4,64'h1da1c8cedc0a82b1,64'h425dc905dd0b407c,64'h5a912f4c44e9ea2f,
64'h6535171c512866cf,64'h789cc293d8dd1a0a,64'h879db5e024bc2928,64'h07fffffffffff800,
64'hfc3f338e2e1be3e1,64'h26872e386bba19e7,64'h1518f92885e5c903,64'h4086b22262f70758,
64'h72a89641095e5008,64'hadf8fb90ab8d79bc,64'hd395a5ae65fc714b,64'h7d17eac4df70590d,
64'h8fad933eddd29733,64'hac7dfbdd8929959e,64'h3a36d11d60e31cc5,64'h9428f55543e67bab,
64'hfbb4631ceff22eb2,64'he6e62d7fdd6029b6,64'h9bfcda44fc5dd883,64'h0b9016d6b8c3f082,
64'hb63d9dbd712b6817,64'h71e22c5fb4cd7de1,64'h9cc738100790eeac,64'h7eed9cffcab60a64,
64'h7f41d0cd8235564c,64'h91d5de15c8589dd1,64'hf408e8f386f8367c,64'hc26e0b997ad762f0,
64'hc3d29b52cdaef7f8,64'h7712092d45a443da,64'h0a4225683671b7d8,64'h3a956717ac822bd5,
64'h1760e239a7ce938c,64'h91911f54f937fdd4,64'hb6f99b31fd512b23,64'hffdfffff00200001
};
  //------------------------
  // 1024
  //------------------------
  localparam [2*1024-1:0][63:0] NTT_GF64_BWD_WDIV_N1024_PHI_L = {
64'h061e96455f799f0a,64'h518f6817aa1c313d,64'hf080d371f8e2b141,64'habf210fbace5182e,
64'h2d7fd707ec6c09cb,64'h428e6beb188ca2c6,64'h7d95bb07123ec141,64'hb4b0b7b3a810dd79,
64'hb55cc38ebf1e85df,64'hd702ff65e35e274a,64'h090e87c90457bc57,64'hf496a73b2d4f9244,
64'hda1c8ceec0a82b0f,64'ha912f4c94e9ea2eb,64'h89cc29448dd1a099,64'h7fffffffffff8000,
64'h6872e388bba19e6e,64'h086b222a2f70757c,64'hdf8fb914b8d79bb6,64'hd17eac54f70590c9,
64'hc7dfbde2929959d6,64'h428f555d3e67baa7,64'h6e62d80bd6029b52,64'hb9016d6b8c3f0820,
64'h1e22c6024cd7de09,64'heed9d003ab60a639,64'h1d5de1658589dd07,64'h26e0b9a3ad762ef4,
64'h712092db5a443d99,64'ha956717dc822bd4d,64'h1911f558937fdd37,64'hfdffffff02000001,
64'h30f4b22afbccf850,64'h8c7b40bf50e189e6,64'h84069b96c7158a01,64'h5f9087e26728c16b,
64'h6bfeb84063604e57,64'h14735f5ac465162e,64'hecadd83b91f60a05,64'ha585bda24086ebc3,
64'haae61c7af8f42ef3,64'hb817fb351af13a4a,64'h48743e4822bde2b8,64'ha4b539e06a7c9219,
64'hd0e4677c05415872,64'h4897a64f74f51753,64'h4e614a286e8d04c4,64'h00000003fffbfffc,
64'h43971c48dd0cf36d,64'h435911517b83abe0,64'hfc7dc8abc6bcddaa,64'h8bf562adb82c8642,
64'h3efdef1a94caceaa,64'h147aaaebf33dd536,64'h7316c061b014da8d,64'hc80b6b6161f840fb,
64'hf116301266bef048,64'h76ce80245b0531c1,64'heaef0b2c2c4ee838,64'h3705cd1e6bb1779f,
64'h890496ddd221ecc5,64'h4ab38bf34115ea63,64'hc88faac49bfee9b8,64'hefffffff10000001,
64'h87a59158de67c27f,64'h63da05fe870c4f2c,64'h2034dcba38ac5004,64'hfc843f1539460b56,
64'h5ff5c2061b0272b5,64'ha39afad62328b170,64'h656ec1e38fb05021,64'h2c2ded1704375e13,
64'h5730e3dcc7a17793,64'hc0bfd9add789d24b,64'h43a1f24315ef15be,64'h25a9cf0853e490c3,
64'h87233be62a0ac38a,64'h44bd327da7a8ba96,64'h730a51457468261e,64'h0000001fffdfffe0,
64'h1cb8e248e8679b66,64'h1ac88a8ddc1d5efe,64'he3ee456535e6ed49,64'h5fab1571c164320c,
64'hf7ef78d5a656754f,64'ha3d5575f99eea9b0,64'h98b6031080a6d465,64'h405b5b110fc207d2,
64'h88b1809a35f78239,64'hb6740125d8298e05,64'h57785968627741b9,64'hb82e68f45d8bbcf7,
64'h4824b6f2910f6624,64'h559c5f9c08af5316,64'h447d562adff74dba,64'h7fffffff80000001,
64'h3d2c8acaf33e13f4,64'h1ed02ff73862795d,64'h01a6e5d2c562801f,64'he421f8b0ca305aa9,
64'hffae1032d81395a6,64'h1cd7d6b619458b7b,64'h2b760f1f7d828105,64'h616f68b921baf097,
64'hb9871ee83d0bbc96,64'h05fecd74bc4e9252,64'h1d0f921aaf78adee,64'h2d4e78439f248617,
64'h3919df3550561c4c,64'h25e993ef3d45d4ae,64'h98528a2ea34130ed,64'h000000fffeffff00,
64'he5c71247433cdb30,64'hd644546ee0eaf7f0,64'h1f722b30af376a41,64'hfd58ab900b21905e,
64'hbf7bc6b432b3aa71,64'h1eaabb01cf754d7b,64'hc5b018880536a324,64'h02dad88a7e103e8e,
64'h458c04d5afbc11c4,64'hb3a00933c14c7023,64'hbbc2cb4513ba0dc6,64'hc17347a7ec5de7b3,
64'h4125b796887b311e,64'hace2fce2457a98ae,64'h23eab158ffba6dce,64'h0000000000000004,
64'he964565899f09f9f,64'hf6817fb9c313cae8,64'h0d372e962b1400f8,64'h210fc58d5182d541,
64'hfd70819dc09cad29,64'he6beb5b0ca2c5bd8,64'h5bb078fcec140827,64'h0b7b45cc0dd784b5,
64'hcc38f746e85de4ab,64'h2ff66ba5e2749290,64'he87c90d57bc56f70,64'h6a73c21df92430b7,
64'hc8cef9ab82b0e25f,64'h2f4c9f7aea2ea56f,64'hc29451791a098764,64'h000007fff7fff800,
64'h2e38924119e6d979,64'hb222a37d0757bf7a,64'hfb91598579bb5208,64'heac55c87590c82e9,
64'hfbde35a6959d5383,64'hf555d80e7baa6bd8,64'h2d80c44629b5191a,64'h16d6c453f081f470,
64'h2c6026af7de08e1e,64'h9d0049a30a638113,64'hde165a2d9dd06e2b,64'h0b9a3d4562ef3d92,
64'h092dbcb643d988ee,64'h6717e7172bd4c56b,64'h1f558ac8fdd36e6f,64'h0000000000000020,
64'h4b22b2cbcf84fcf1,64'hb40bfdd5189e5739,64'h69b974b158a007c0,64'h087e2c6b8c16aa07,
64'heb840cf504e56941,64'h35f5ad8d5162deb9,64'hdd83c7e960a04136,64'h5bda2e606ebc25a8,
64'h61c7ba3d42ef2552,64'h7fb35d3013a4947f,64'h43e486b2de2b7b79,64'h539e10f2c92185b5,
64'h4677cd62158712f2,64'h7a64fbd851752b77,64'h14a28bced04c3b1a,64'h00003fffbfffc000,
64'h71c49209cf36cbc7,64'h91151bed3abdfbcb,64'hdc8acc32cdda9039,64'h562ae441c8641741,
64'hdef1ad3bacea9c11,64'haaaec07add535eb9,64'h6c0622324da8c8cf,64'hb6b6229f840fa380,
64'h6301357cef0470ef,64'he8024d1c531c0894,64'hf0b2d172ee837152,64'h5cd1ea2b1779ec90,
64'h496de5b21ecc4770,64'h38bf38bc5ea62b55,64'hfaac5647ee9b7378,64'h0000000000000100,
64'h591596607c27e786,64'ha05feeadc4f2b9c3,64'h4dcba58dc5003dfd,64'h43f1635c60b55038,
64'h5c2067af272b4a01,64'hafad6c6b8b16f5c7,64'hec1e3f51050209aa,64'hded1730575e12d3e,
64'h0e3dd1ed17792a8d,64'hfd9ae9839d24a3f5,64'h1f243598f15bdbc6,64'h9cf08798490c2da6,
64'h33be6b12ac38978e,64'hd327dec58ba95bb5,64'ha5145e768261d8d0,64'h0001fffdfffe0000,
64'h8e24905179b65e35,64'h88a8df6dd5efde54,64'he456619c6ed481c2,64'hb15722104320ba06,
64'hf78d69e36754e082,64'h557603dbea9af5c3,64'h603111956d464675,64'hb5b11501207d1bfb,
64'h1809abea78238775,64'h401268e998e04499,64'h85968b9e741b8a89,64'he68f515abbcf647e,
64'h4b6f2d92f6623b7e,64'hc5f9c5e3f5315aa7,64'hd562b24674db9bb9,64'h0000000000000800,
64'hc8acb305e13f3c2e,64'h02ff75732795ce13,64'h6e5d2c702801efe6,64'h1f8b1ae505aa81be,
64'he1033d7b395a5006,64'h7d6b636158b7ae33,64'h60f1fa8f28104d49,64'hf68b9831af0969ea,
64'h71ee8f68bbc95468,64'hecd74c23e9251fa1,64'hf921acc78adede30,64'he7843cc648616d2c,
64'h9df3589661c4bc6f,64'h993ef6325d4adda2,64'h28a2f3b9130ec67b,64'h000fffeffff00000,
64'h7124828fcdb2f1a4,64'h4546fb72af7ef29c,64'h22b30cea76a40e09,64'h8ab910871905d02b,
64'hbc6b4f223aa70409,64'habb01ee154d7ae16,64'h01888cae6a3233a5,64'had88a80e03e8dfd3,
64'hc04d5f53c11c3ba8,64'h0093474ec70224c6,64'h2cb45cf7a0dc5444,64'h347a8adcde7b23e9,
64'h5b796c99b311dbee,64'h2fce2f25a98ad532,64'hab159239a6dcddc2,64'h0000000000004000,
64'h4565983509f9e16a,64'h17fbab993cae7098,64'h72e96384400f7f2d,64'hfc58d7282d540df0,
64'h0819ebe0cad28029,64'heb5b1b0dc5bd7195,64'h078fd47c40826a45,64'hb45cc194784b4f49,
64'h8f747b48de4aa33d,64'h66ba61264928fd01,64'hc90d664356f6f179,64'h3c21e639430b6959,
64'hef9ac4b70e25e374,64'hc9f7b196ea56ed0c,64'h45179dc9987633d7,64'h007fff7fff800000,
64'h892414816d978d1d,64'h2a37db977bf794de,64'h15986754b5207047,64'h55c8843cc82e8154,
64'he35a7916d5382043,64'h5d80f70fa6bd70ab,64'h0c44657351919d28,64'h6c4540751f46fe93,
64'h026afaa408e1dd3a,64'h049a3a7638112630,64'h65a2e7be06e2a21f,64'ha3d456e7f3d91f47,
64'hdbcb64cf988edf6e,64'h7e71792e4c56a98f,64'h58ac91d236e6ee0b,64'h0000000000020000,
64'h2b2cc1aa4fcf0b4e,64'hbfdd5cc9e57384c0,64'h974b1c25007bf965,64'he2c6b9486aa06f79,
64'h40cf5f0656940148,64'h5ad8d8752deb8ca1,64'h3c7ea3e204135228,64'ha2e60ca8c25a7a43,
64'h7ba3da4af25519e4,64'h35d309354947e805,64'h486b3220b7b78bc2,64'he10f31cb185b4ac7,
64'h7cd625bf712f1b99,64'h4fbd8cbd52b7685a,64'h28bcee4ec3b19eb6,64'h03fffbfffc000000,
64'h4920a40f6cbc68e4,64'h51bedcbcdfbca6ef,64'hacc33aa5a9038238,64'hae4421e841740a9e,
64'h1ad3c8bda9c10211,64'hec07b87f35eb8556,64'h62232b9a8c8ce940,64'h622a03abfa37f495,
64'h1357d520470ee9d0,64'h24d1d3b1c0893180,64'h2d173df3371510f5,64'h1ea2b7449ec8fa33,
64'hde5b2682c476fb6a,64'hf38bc97562b54c75,64'hc5648e93b7377056,64'h0000000000100000,
64'h59660d537e785a6f,64'hfeeae6542b9c25fb,64'hba58e12c03dfcb24,64'h1635ca4a55037bc1,
64'h067af834b4a00a3e,64'hd6c6c3ab6f5c6506,64'he3f51f11209a913f,64'h1730654b12d3d213,
64'hdd1ed25a92a8cf1d,64'hae9849ab4a3f4027,64'h43599107bdbc5e0e,64'h08798e5fc2da5631,
64'he6b12dfe8978dcc5,64'h7dec65ec95bb42ce,64'h45e772771d8cf5af,64'h1fffdfffe0000000,
64'h4905207d65e3471e,64'h8df6e5e8fde53776,64'h6619d532481c11bb,64'h72210f470ba054eb,
64'hd69e45ed4e081088,64'h603dc400af5c2aa9,64'h11195cd7646749fd,64'h11501d62d1bfa4a5,
64'h9abea90238774e80,64'h268e9d8f04498bff,64'h68b9ef9ab8a887a7,64'hf515ba24f647d198,
64'hf2d9341c23b7db4a,64'h9c5e4bb215aa63a1,64'h2b2474a3b9bb82aa,64'h0000000000800000,
64'hcb306a9df3c2d376,64'hf75732a85ce12fd1,64'hd2c709651efe591b,64'hb1ae5252a81bde08,
64'h33d7c1a5a50051f0,64'hb6361d617ae3282a,64'h1fa8f89004d489f1,64'hb9832a58969e9098,
64'he8f692da954678e2,64'h74c24d5f51fa0133,64'h1acc883fede2f06e,64'h43cc72fe16d2b188,
64'h35896ffb4bc6e621,64'hef632f67adda166d,64'h2f3b93baec67ad76,64'hfffeffff00000000,
64'h482903ed2f1a38ee,64'h6fb72f4bef29bbac,64'h30cea99540e08dd5,64'h91087a3b5d02a755,
64'hb4f22f707040843a,64'h01ee20087ae15545,64'h88cae6bb233a4fe8,64'h8a80eb168dfd2528,
64'hd5f54815c3ba73fc,64'h3474ec79224c5ff7,64'h45cf7cd8c5443d35,64'ha8add12eb23e8cb9,
64'h96c9a0e81dbeda49,64'he2f25d94ad531d04,64'h5923a51ecddc154f,64'h0000000004000000,
64'h598354f59e169baa,64'hbab99549e7097e81,64'h96384b2ef7f2c8d2,64'h8d72929a40def03b,
64'h9ebe0d2e28028f7f,64'hb1b0eb10d719414b,64'hfd47c48026a44f88,64'hcc1952c9b4f484bb,
64'h47b496dbaa33c709,64'ha6126afd8fd00995,64'hd66441ff6f178370,64'h1e6397f2b6958c3e,
64'hac4b7fdb5e373107,64'h7b197b446ed0b361,64'h79dc9dd8633d6baf,64'hfff7fffefffffff9,
64'h41481f6b78d1c76e,64'h7db97a62794ddd5d,64'h86754cab07046ea7,64'h8843d1dee8153aa4,
64'ha7917b88820421cb,64'h0f710043d70aaa28,64'h465735dd19d27f3c,64'h540758b86fe9293c,
64'hafaa40b41dd39fda,64'ha3a763ca1262ffb7,64'h2e7be6c82a21e9a6,64'h456e897a91f465c3,
64'hb64d0744edf6d244,64'h1792ecac6a98e819,64'hc91d28f86ee0aa76,64'h0000000020000000,
64'hcc1aa7aef0b4dd4e,64'hd5ccaa54384bf403,64'hb1c2597bbf96468c,64'h6b9494d606f781d4,
64'hf5f0697540147bf4,64'h8d87588bb8ca0a53,64'hea3e240835227c39,64'h60ca9653a7a425d2,
64'h3da4b6df519e3846,64'h309357f17e804ca3,64'hb322100178bc1b7a,64'hf31cbf95b4ac61f0,
64'h625bfedff1b98833,64'hd8cbda2676859b05,64'hcee4eec619eb5d75,64'hffbffffeffffffc1,
64'h0a40fb5dc68e3b6e,64'hedcbd316ca6eeae5,64'h33aa655c38237534,64'h421e8efb40a9d51c,
64'h3c8bdc4910210e53,64'h7b88021eb8555140,64'h32b9aeeace93f9de,64'ha03ac5c57f4949de,
64'h7d5205a5ee9cfecb,64'h1d3b1e559317fdb3,64'h73df3642510f4d2f,64'h2b744bd68fa32e16,
64'hb2683a2c6fb6921b,64'hbc97656354c740c8,64'h48e947c9770553aa,64'h0000000100000000,
64'h60d53d7d85a6ea6a,64'hae6552a7c25fa012,64'h8e12cbe2fcb2345b,64'h5ca4a6b337bc0e9d,
64'haf834bb100a3df99,64'h6c3ac461c6505294,64'h51f12048a913e1c1,64'h0654b2a03d212e8d,
64'hed25b6fb8cf1c22f,64'h849abf8cf4026517,64'h99108010c5e0dbcb,64'h98e5fcb4a5630f79,
64'h12dff7028dcc4195,64'hc65ed139b42cd822,64'h77277636cf5aeba2,64'hfdfffffefffffe01,
64'h5207daee3471db70,64'h6e5e98bd53775721,64'h9d532ae2c11ba99f,64'h10f477dc054ea8de,
64'he45ee24981087297,64'hdc4010f8c2aa89fd,64'h95cd7757749fceef,64'h01d62e30fa4a4eeb,
64'hea902d3274e7f655,64'he9d8f2ac98bfed98,64'h9ef9b215887a6975,64'h5ba25eb57d1970af,
64'h9341d1687db490d3,64'he4bb2b1fa63a063b,64'h474a3e4db82a9d4e,64'h0000000800000000,
64'h06a9ebef2d37534d,64'h732a954312fd008b,64'h70965f1be591a2d4,64'he525359bbde074e6,
64'h7c1a5d8d051efcc3,64'h61d623113282949d,64'h8f890247489f0e06,64'h32a59501e9097468,
64'h692db7e3678e1171,64'h24d5fc6ba01328b4,64'hc884008a2f06de54,64'hc72fe5a92b187bc4,
64'h96ffb8146e620ca8,64'h32f689d3a166c10a,64'hb93bb1b97ad75d0d,64'heffffffefffff001,
64'h903ed773a38edb7e,64'h72f4c5ed9bbab905,64'hea99571a08dd4cf4,64'h87a3bee02a7546f0,
64'h22f71253084394b1,64'he20087cc15544fe2,64'hae6bbabfa4fe7774,64'h0eb17187d2527758,
64'h5481699aa73fb2a1,64'h4ec7956bc5ff6cb9,64'hf7cd90b043d34ba4,64'hdd12f5ade8cb8576,
64'h9a0e8b47eda48694,64'h25d9590431d031d1,64'h3a51f26fc154ea6e,64'h0000004000000000,
64'h354f5f7969ba9a68,64'h9954aa1b97e80455,64'h84b2f8e22c8d169d,64'h2929ace4ef03a729,
64'he0d2ec6b28f7e615,64'h0eb1188c9414a4e5,64'h7c48123e44f8702c,64'h952ca810484ba33f,
64'h496dbf1e3c708b85,64'h26afe35e0099459f,64'h442004577836f29a,64'h397f2d4f58c3de1a,
64'hb7fdc0a77310653c,64'h97b44e9e0b36084f,64'hc9dd8dd0d6bae863,64'h7ffffffeffff8001,
64'h81f6bba11c76dbec,64'h97a62f6fddd5c825,64'h54cab8d746ea6799,64'h3d1df70553aa377c,
64'h17b89299421ca587,64'h10043e67aaa27f09,64'h735dd60227f3bb9b,64'h758b8c3e9293bac0,
64'ha40b4cd739fd9506,64'h763cab602ffb65c6,64'hbe6c85891e9a5d19,64'he897ad75465c2baa,
64'hd0745a436d24349c,64'h2ecac8228e818e87,64'hd28f937f0aa7536f,64'h0000020000000000,
64'haa7afbcc4dd4d33f,64'hcaa550e0bf4022a4,64'h2597c7156468b4e4,64'h494d6728781d3947,
64'h0697636047bf30a1,64'h7588c464a0a52728,64'he24091f527c3815d,64'ha9654086425d19f4,
64'h4b6df8f3e3845c26,64'h357f1af104ca2cf7,64'h210022bdc1b794ce,64'hcbf96a7bc61ef0cf,
64'hbfee0540988329db,64'hbda274f459b04274,64'h4eec6e8cb5d74312,64'hfffffffafffc0005,
64'h0fb5dd0ce3b6df5c,64'hbd317b82eeae4124,64'ha655c6bc37533cc6,64'he8efb82b9d51bbdf,
64'hbdc494ca10e52c38,64'h8021f33d5513f848,64'h9aeeb0143f9ddcd5,64'hac5c61f7949dd5fd,
64'h205a66becfeca82b,64'hb1e55b047fdb2e2d,64'hf3642c4df4d2e8c3,64'h44bd6bb132e15d49,
64'h83a2d2216921a4da,64'h76564115740c7437,64'h947c9bfe553a9b72,64'h0000100000000000,
64'h53d7de676ea699f3,64'h552a870bfa01151a,64'h2cbe38ac2345a71f,64'h4a6b3945c0e9ca36,
64'h34bb1b023df98508,64'hac4623280529393d,64'h12048fb03e1c0ae1,64'h4b2a043712e8cf9b,
64'h5b6fc7a11c22e12e,64'habf8d789265167b7,64'h080115ef0dbca66f,64'h5fcb53e430f78672,
64'hff702a09c4194ed3,64'hed13a7a7cd82139b,64'h77637467aeba188e,64'hffffffdeffe00021,
64'h7daee8671db6fae0,64'he98bdc1c7572091b,64'h32ae35e6ba99e62b,64'h477dc163ea8ddef1,
64'hee24a655872961bb,64'h010f99eea89fc23c,64'hd77580a5fceee6a4,64'h62e30fc1a4eeafe3,
64'h02d335f77f654157,64'h8f2ad828fed97163,64'h9b216276a6974611,64'h25eb5d8b970aea46,
64'h1d16910f490d26cc,64'hb2b208aea063a1b5,64'ha3e4dff6a9d4db8c,64'h0000800000000000,
64'h9ebef33d7534cf96,64'ha9543861d008a8ce,64'h65f1c5621a2d38f7,64'h5359ca30074e51ae,
64'ha5d8d812efcc283f,64'h623119452949c9e3,64'h90247d81f0e05708,64'h595021ba97467cd6,
64'hdb7e3d0ae117096e,64'h5fc6bc4e328b3db3,64'h4008af786de53378,64'hfe5a9f2387bc338e,
64'hfb81505520ca7691,64'h689d3d456c109cd1,64'hbb1ba34075d0c46d,64'hfffffefeff000101,
64'hed77433bedb7d6fd,64'h4c5ee0eaab9048d1,64'h9571af36d4cf3157,64'h3bee0b21546ef786,
64'h712532b3394b0dd1,64'h087ccf7544fe11e0,64'hbbac0535e777351a,64'h17187e1027757f15,
64'h1699afbbfb2a0ab8,64'h7956c14bf6cb8b14,64'hd90b13b934ba3084,64'h2f5aec5db857522f,
64'he8b4887a48693660,64'h9590457a031d0da3,64'h1f26ffba4ea6dc5b,64'h0004000000000000,
64'hf5f799efa9a67cac,64'h4aa1c3138045466b,64'h2f8e2b13d169c7b5,64'h9ace51823a728d6e,
64'h2ec6c09c7e6141f3,64'h1188ca2c4a4e4f15,64'h8123ec138702b83c,64'hca810dd6ba33e6ae,
64'hdbf1e85d08b84b6a,64'hfe35e2739459ed96,64'h00457bc56f299bbe,64'hf2d4f9233de19c69,
64'hdc0a82b00653b481,64'h44e9ea2e6084e685,64'hd8dd1a08ae862363,64'hfffff7fef8000801,
64'h6bba19e66dbeb7e1,64'h62f707575c824686,64'hab8d79baa6798ab4,64'hdf70590ba377bc2f,
64'h8929959cca586e85,64'h43e67baa27f08f00,64'hdd6029b43bb9a8cb,64'hb8c3f0813babf8a8,
64'hb4cd7ddfd95055c0,64'hcab60a62b65c589d,64'hc8589dcfa5d1841a,64'h7ad762eec2ba9177,
64'h45a443d94349b2f9,64'hac822bd418e86d14,64'hf937fdd27536e2d8,64'h0020000000000000,
64'hafbccf844d33e559,64'h550e189e022a3356,64'h7c71589f8b4e3da7,64'hd6728c15d3946b6c,
64'h763604e4f30a0f97,64'h8c465162527278a8,64'h091f60a03815c1dc,64'h54086ebbd19f356a,
64'hdf8f42ee45c25b4a,64'hf1af13a3a2cf6ca9,64'h022bde2b794cddf0,64'h96a7c920ef0ce341,
64'he0541586329da402,64'h274f517504273426,64'hc6e8d04b74311b12,64'hffffbffec0004001,
64'h5dd0cf366df5bf05,64'h17b83abde412342d,64'h5c6bcdda33cc559b,64'hfb82c8631bbde172,
64'h494cacea52c37424,64'h1f33dd533f8477fe,64'heb014da7ddcd4652,64'hc61f840edd5fc53b,
64'ha66bef03ca82adfb,64'h55b0531bb2e2c4e2,64'h42c4ee832e8c20ca,64'hd6bb177915d48bb5,
64'h2d221ecc1a4d97c6,64'h64115ea5c743689b,64'hc9bfee9aa9b716b9,64'h0100000000000000,
64'h7de67c27699f2ac3,64'ha870c4f211519aae,64'he38ac4ff5a71ed35,64'hb39460b49ca35b5a,
64'hb1b0272a98507cb5,64'h62328b169393c53c,64'h48fb0501c0ae0ee0,64'ha04375e08cf9ab4e,
64'hfc7a17782e12da4a,64'h8d789d24167b6541,64'h115ef15bca66ef80,64'hb53e490b78671a04,
64'h02a0ac3894ed2009,64'h3a7a8ba92139a12f,64'h37468261a188d88a,64'hfffdfffd00020001,
64'hee8679b56fadf826,64'hbdc1d5ef2091a168,64'he35e6ed39e62acd6,64'hdc16431fddef0b89,
64'h4a656754961ba11e,64'hf99eea99fc23bff0,64'h580a6d45ee6a3289,64'h30fc207ceafe29d2,
64'h335f782354156fd3,64'had8298df9716270e,64'h1627741b7461064e,64'hb5d8bbceaea45da2,
64'h6910f661d26cbe2f,64'h208af5313a1b44d5,64'h4dff74db4db8b5c2,64'h0800000000000000,
64'hef33e13e4cf95615,64'h438627958a8cd56b,64'h1c562801d38f69a1,64'h9ca305a9e51adacb,
64'h8d813959c283e5a3,64'h119458b79c9e29dd,64'h47d82810057076fe,64'h021baf0967cd5a6b,
64'he3d0bbc87096d249,64'h6bc4e924b3db2a04,64'h8af78ade53377c00,64'ha9f24860c338d01b,
64'h150561c4a7690048,64'hd3d45d4a09cd0977,64'hba34130e0c46c44f,64'hffefffef00100001,
64'h7433cdb27d6fc129,64'hee0eaf7e048d0b3b,64'h1af376a3f31566a9,64'he0b21904ef785c42,
64'h532b3aa6b0dd08ee,64'hccf754d6e11dff79,64'hc0536a3173519446,64'h87e103e857f14e8f,
64'h9afbc11ba0ab7e97,64'h6c14c701b8b1386b,64'hb13ba0dba3083270,64'haec5de7a7522ed0b,
64'h4887b3119365f175,64'h0457a98ad0da26a7,64'h6ffba6dc6dc5ae0e,64'h4000000000000000,
64'h799f09f967cab0a1,64'h1c313cae5466ab56,64'he2b1400e9c7b4d08,64'he5182d5328d6d654,
64'h6c09cad2141f2d14,64'h8ca2c5bce4f14ee8,64'h3ec140822b83b7ee,64'h10dd784b3e6ad358,
64'h1e85de4a84b69241,64'h5e2749289ed9501d,64'h57bc56f699bbdffc,64'h4f92430b19c680d3,
64'ha82b0e253b480240,64'h9ea2ea564e684bb2,64'hd1a0987562362273,64'hff7fff7f00800001,
64'ha19e6d96eb7e0945,64'h70757bf7246859d1,64'hd79bb51f98ab3548,64'h0590c82e7bc2e209,
64'h9959d53786e8476e,64'h67baa6bd08effbc2,64'h029b51919a8ca22a,64'h3f081f46bf8a7474,
64'hd7de08e1055bf4b4,64'h60a63810c589c355,64'h89dd06e21841937b,64'h762ef3d8a9176853,
64'h443d988e9b2f8ba6,64'h22bd4c5686d13538,64'h7fdd36e66e2d706d,64'h00000001fffffffe,
64'hccf84fce3e558505,64'he189e572a3355ab0,64'h158a007be3da6839,64'h28c16aa046b6b299,
64'h604e5693a0f9689d,64'h65162deb278a773c,64'hf60a04125c1dbf6f,64'h86ebc259f3569ac0,
64'hf42ef25425b49208,64'hf13a4946f6ca80e6,64'hbde2b7b6cddeffde,64'h7c92185ace340696,
64'h4158712eda4011fb,64'hf51752b673425d8c,64'h8d04c3b111b11392,64'hfbfffbff04000001,
64'h0cf36cbc5bf04a23,64'h83abdfbc2342ce85,64'hbcdda902c559aa3a,64'h2c864173de171048,
64'hcacea9c037423b6c,64'h3dd535eb477fde0d,64'h14da8c8cd4651150,64'hf840fa36fc53a39f,
64'hbef0470e2adfa59a,64'h0531c0892c4e1aa5,64'h4ee83714c20c9bd4,64'hb1779ec848bb4295,
64'h21ecc476d97c5d2e,64'h15ea62b53689a9bf,64'hfee9b736716b8365,64'h0000000ffffffff0,
64'h67c27e77f2ac2822,64'h0c4f2b9c19aad579,64'hac5003df1ed341c8,64'h460b550335b594c7,
64'h0272b4a007cb44e5,64'h28b16f5c3c53b9dd,64'hb0502099e0edfb71,64'h375e12d39ab4d5fc,
64'ha17792a82da49039,64'h89d24a3eb6540729,64'hef15bdbb6ef7feeb,64'he490c2d971a034ad,
64'h0ac38978d2008fd6,64'ha8ba95ba9a12ec59,64'h68261d8c8d889c8c,64'hdfffdfff20000001,
64'h679b65e2df825118,64'h1d5efde51a167424,64'he6ed481b2acd51cb,64'h64320b9ff0b8823f,
64'h56754e07ba11db5a,64'heea9af5b3bfef067,64'ha6d46466a3288a80,64'hc207d1bee29d1cf1,
64'hf782387656fd2ccb,64'h298e04496270d528,64'h7741b8a81064de9e,64'h8bbcf64745da14a3,
64'h0f6623b7cbe2e96f,64'haf5315a9b44d4df8,64'hf74db9ba8b5c1b21,64'h0000007fffffff80,
64'h3e13f3c29561410d,64'h62795ce0cd56abc8,64'h62801efdf69a0e3b,64'h305aa81badaca636,
64'h1395a5003e5a2728,64'h458b7ae2e29dcee7,64'h828104d4076fdb83,64'hbaf0969dd5a6afdf,
64'h0bbc95466d2481c3,64'h4e9251f9b2a03944,64'h78adede277bff751,64'h248616d28d01a561,
64'h561c4bc690047eb0,64'h45d4add9d09762c3,64'h4130ec676c44e45d,64'hfffeffff00000002,
64'h3cdb2f19fc1288bd,64'heaf7ef28d0b3a120,64'h376a40e0566a8e51,64'h21905d0285c411f5,
64'hb3aa703fd08edace,64'h754d7ae0dff78331,64'h36a3233a194453fb,64'h103e8dfd14e8e782,
64'hbc11c3b9b7e96651,64'h4c70224c1386a93f,64'hba0dc5438326f4ed,64'h5de7b23e2ed0a514,
64'h7b311dbe5f174b78,64'h7a98ad52a26a6fbb,64'hba6dcddb5ae0d901,64'h000003fffffffc00,
64'hf09f9e15ab0a0867,64'h13cae7096ab55e3d,64'h1400f7f2b4d071d5,64'h82d540de6d6531af,
64'h9cad2801f2d13940,64'h2c5bd71914ee7736,64'h140826a43b7edc14,64'hd784b4f3ad357ef3,
64'h5de4aa3369240e18,64'h74928fcf9501ca1e,64'hc56f6f16bdffba85,64'h2430b695680d2b07,
64'hb0e25e368023f57e,64'h2ea56ed084bb1616,64'h0987633d622722e6,64'hfff7ffff00000009,
64'he6d978d0e09445e7,64'h57bf794d859d08f9,64'hbb520703b3547287,64'h0c82e8152e208fa7,
64'h9d5382038476d66b,64'haa6bd709ffbc1985,64'hb51919d1ca229fd7,64'h81f46fe8a7473c10,
64'he08e1dd2bf4b3283,64'h638112629c3549f6,64'hd06e2a211937a763,64'hef3d91f37685289e,
64'hd988edf5f8ba5bbd,64'hd4c56a9813537dd5,64'hd36e6edfd706c803,64'h00001fffffffe000,
64'h84fcf0b458504331,64'h9e57384b55aaf1e8,64'ha007bf95a6838ea8,64'h16aa06f76b298d74,
64'he56940139689c9fc,64'h62deb8c9a773b9af,64'ha0413521dbf6e0a0,64'hbc25a7a369abf792,
64'hef25519d492070be,64'ha4947e7fa80e50ed,64'h2b7b78bbeffdd422,64'h2185b4ac40695837,
64'h8712f1b9011fabeb,64'h752b768525d8b0af,64'h4c3b19eb11391730,64'hffbfffff00000041,
64'h36cbc68e04a22f31,64'hbdfbca6e2ce847c6,64'hda9038229aa39433,64'h641740a971047d38,
64'hea9c102023b6b354,64'h535eb854fde0cc23,64'ha8c8ce935114feb3,64'h0fa37f493a39e07c,
64'h0470ee9cfa599411,64'h1c089317e1aa4fad,64'h8371510ec9bd3b12,64'h79ec8fa2b42944e9,
64'hcc476fb5c5d2dde2,64'ha62b54c69a9beea2,64'h9b737704b8364012,64'h0000ffffffff0000,
64'h27e785a6c2821984,64'hf2b9c25ead578f3c,64'h003dfcb2341c753b,64'hb55037bb594c6ba0,
64'h2b4a00a3b44e4fd9,64'h16f5c6503b9dcd75,64'h0209a913dfb704fb,64'he12d3d204d5fbc8b,
64'h792a8cf1490385e9,64'h24a3f40240728763,64'h5bdbc5e07feea10f,64'h0c2da563034ac1b7,
64'h38978dcc08fd5f54,64'ha95bb42c2ec58575,64'h61d8cf5a89c8b97e,64'hfdffffff00000201,
64'hb65e347125117987,64'hefde537667423e2b,64'hd481c11ad51ca192,64'h20ba054e8823e9bd,
64'h54e081081db59a99,64'h9af5c2a9ef066116,64'h4646749f88a7f593,64'h7d1bfa49d1cf03e0,
64'h238774e7d2cca088,64'he04498bf0d527d68,64'h1b8a887a4de9d88c,64'hcf647d18a14a2745,
64'h623b7db42e96ef0a,64'h315aa639d4df750b,64'hdb9bb829c1b2008c,64'h0007fffffff80000,
64'h3f3c2d371410cc1f,64'h95ce12fc6abc79d9,64'h01efe591a0e3a9d8,64'haa81bddfca635cfb,
64'h5a50051ea2727ec7,64'hb7ae3281dcee6ba8,64'h104d489efdb827d8,64'h0969e9096afde451,
64'hc954678d481c2f45,64'h251fa01303943b17,64'hdede2f05ff750876,64'h616d2b181a560db8,
64'hc4bc6e6147eafa9f,64'h4adda166762c2ba3,64'h0ec67ad74e45cbed,64'hefffffff00001001,
64'hb2f1a38e288bcc33,64'h7ef29bba3a11f151,64'ha40e08dca8e50c8a,64'h05d02a75411f4de7,
64'ha7040842edacd4c6,64'hd7ae1553783308ac,64'h3233a4fe453fac96,64'he8dfd2518e781efd,
64'h1c3ba73f9665043f,64'h0224c5ff6a93eb39,64'hdc5443d26f4ec460,64'h7b23e8cb0a513a22,
64'h11dbeda474b7784d,64'h8ad531cfa6fba857,64'hdcddc1540d90045a,64'h003fffffffc00000,
64'hf9e169b9a08660f7,64'hae7097e755e3cec4,64'h0f7f2c8d071d4ec0,64'h540def03531ae7d3,
64'hd28028f71393f636,64'hbd719413e7735d3b,64'h826a44f7edc13ec0,64'h4b4f484b57ef2288,
64'h4aa33c7040e17a22,64'h28fd00991ca1d8b7,64'hf6f17835fba843aa,64'h0b6958c3d2b06dbd,
64'h25e373103f57d4f2,64'h56ed0b35b1615d16,64'h7633d6ba722e5f68,64'h7fffffff00008001,
64'h978d1c76445e6193,64'hf794ddd4d08f8a85,64'h207046ea4728644b,64'h2e8153aa08fa6f38,
64'h3820421c6d66a62b,64'hbd70aaa1c198455a,64'h919d27f329fd64af,64'h46fe929373c0f7e1,
64'he1dd39fcb32821f8,64'h11262ffb549f59c8,64'he2a21e997a7622fa,64'hd91f465b5289d10d,
64'h8edf6d23a5bbc268,64'h56a98e8137dd42b4,64'he6ee0aa66c8022ca,64'h01fffffffe000000,
64'hcf0b4dd4043307b1,64'h7384bf3faf1e761b,64'h7bf9646838ea7600,64'ha06f781c98d73e96,
64'h940147be9c9fb1aa,64'heb8ca0a43b9ae9d3,64'h135227c36e09f5fc,64'h5a7a425cbf79143e,
64'h5519e384070bd10e,64'h47e804c9e50ec5b7,64'hb78bc1b6dd421d49,64'h5b4ac61e95836de8,
64'h2f1b9882fabea78f,64'hb76859af8b0ae8ae,64'hb19eb5d69172fb3d,64'hfffffffb00040005,
64'hbc68e3b622f30c94,64'hbca6eead847c5421,64'h0382375339432257,64'h740a9d5147d379bf,
64'hc10210e46b353157,64'heb8555130cc22acb,64'h8ce93f9d4feb2574,64'h37f4949d9e07bf06,
64'h0ee9cfec99410fb9,64'h89317fdaa4face40,64'h1510f4d2d3b117c9,64'hc8fa32e0944e8862,
64'h76fb69212dde133c,64'hb54c740bbeea159e,64'h3770553a64011649,64'h0ffffffff0000000,
64'h785a6ea621983d82,64'h9c25fa0078f3b0d5,64'hdfcb2344c753affd,64'h037bc0e9c6b9f4ab,
64'ha00a3df8e4fd8d4c,64'h5c650528dcd74e91,64'h9a913e1b704fafe0,64'hd3d212e7fbc8a1ee,
64'ha8cf1c22385e886e,64'h3f40265128762db6,64'hbc5e0dbbea10ea43,64'hda5630f6ac1b6f3e,
64'h78dcc418d5f53c77,64'hbb42cd815857456b,64'h8cf5aeb98b97d9e3,64'hffffffdf00200021,
64'he3471db61798649b,64'he537757123e2a103,64'h1c11ba99ca1912b8,64'ha054ea8d3e9bcdf5,
64'h0810872959a98ab2,64'h5c2aa89f66115651,64'h6749fcee7f592b9c,64'hbfa4a4edf03df82f,
64'h774e7f64ca087dc8,64'h498bfed927d671fc,64'ha887a6969d88be48,64'h47d1970aa274430a,
64'hb7db490c6ef099dd,64'haa63a062f750aceb,64'hbb82a9d42008b247,64'h7fffffff80000000,
64'hc2d375340cc1ec0d,64'he12fd007c79d86a4,64'hfe591a2c3a9d7fe2,64'h1bde074e35cfa558,
64'h0051efcc27ec6a5b,64'he3282948e6ba7486,64'hd489f0df827d7efc,64'h9e909745de450f6a,
64'h4678e116c2f4436b,64'hfa01328a43b16daf,64'he2f06de450875213,64'hd2b187bb60db79ea,
64'hc6e620c9afa9e3b5,64'hda166c0fc2ba2b53,64'h67ad75d05cbecf14,64'hfffffeff01000101,
64'h1a38edb7bcc324d1,64'h29bbab901f150811,64'he08dd4ce50c895c0,64'h02a7546ef4de6fa3,
64'h4084394acd4c5590,64'he15544fd308ab286,64'h3a4fe776fac95cdd,64'hfd25277481efc173,
64'hba73fb295043ee3d,64'h4c5ff6cb3eb38fde,64'h443d34b9ec45f23b,64'h3e8cb85713a2184e,
64'hbeda48687784cee3,64'h531d031cba856753,64'hdc154ea600459233,64'hfffffffefffffffd,
64'h169ba9a6660f6062,64'h097e80453cec3519,64'hf2c8d168d4ebff09,64'hdef03a71ae7d2ac0,
64'h028f7e613f6352d8,64'h19414a4e35d3a429,64'ha44f870213ebf7da,64'hf484ba32f2287b4c,
64'h33c708b817a21b56,64'hd00994591d8b6d71,64'h17836f29843a9091,64'h958c3de106dbcf4a,
64'h373106537d4f1da2,64'hd0b3608415d15a92,64'h3d6bae85e5f6789d,64'hfffff7ff08000801,
64'hd1c76dbde6192688,64'h4ddd5c81f8a84087,64'h046ea6798644adf9,64'h153aa377a6f37d18,
64'h0421ca586a62ac7e,64'h0aaa27f084559429,64'hd27f3bb8d64ae6e7,64'he9293bab0f7e0b91,
64'hd39fd94f821f71e3,64'h62ffb65bf59c7eee,64'h21e9a5d1622f91d6,64'hf465c2b99d10c26f,
64'hf6d24348bc267713,64'h98e818e7d42b3a96,64'he0aa7536022c9192,64'hfffffffeffffffe1,
64'hb4dd4d33307b0310,64'h4bf40229e761a8c8,64'h96468b4da75ff841,64'hf781d39373e955fa,
64'h147bf309fb1a96c0,64'hca0a5271ae9d2148,64'h227c38159f5fbecb,64'ha425d19e9143da59,
64'h9e3845c1bd10daaf,64'h804ca2ceec5b6b82,64'hbc1b794c21d48488,64'hac61ef0c36de7a4c,
64'hb988329cea78ed0f,64'h859b0426ae8ad48a,64'heb5d74302fb3c4e7,64'hffffbfff40004001,
64'h8e3b6df530c9343a,64'h6eeae411c5420436,64'h237533cc32256fc8,64'ha9d51bbd379be8c0,
64'h210e52c3531563f0,64'h55513f8422aca148,64'h93f9ddccb2573732,64'h4949dd5f7bf05c81,
64'h9cfeca8210fb8f12,64'h17fdb2e2ace3f76d,64'h0f4d2e8c117c8eaf,64'ha32e15d3e8861371,
64'hb6921a4ce133b891,64'hc740c742a159d4ac,64'h0553a9b711648c89,64'hfffffffeffffff01,
64'ha6ea699e83d8187b,64'h5fa011513b0d463e,64'hb2345a713affc204,64'hbc0e9ca29f4aafc9,
64'ha3df984fd8d4b600,64'h5052939374e90a3a,64'h13e1c0adfafdf657,64'h212e8cf98a1ed2c3,
64'hf1c22e11e886d574,64'h0265167b62db5c0c,64'he0dbca660ea4243b,64'h630f7866b6f3d25b,
64'hcc4194ec53c76873,64'h2cd821397456a44c,64'h5aeba1887d9e2731,64'hfffe000100020001,
64'h71db6fad8649a1cc,64'h775720912a1021ad,64'h1ba99e62912b7e3f,64'h4ea8ddeebcdf45fb,
64'h0872961b98ab1f7f,64'haa89fc2315650a3e,64'h9fceee6992b9b98c,64'h4a4eeafddf82e406,
64'he7f6541487dc788c,64'hbfed9715671fbb68,64'h7a6974608be47578,64'h1970aea444309b83,
64'hb490d26c099dc483,64'h3a063a1b0acea55a,64'h2a9d4db88b246448,64'hfffffffefffff801,
64'h37534cf91ec0c3d3,64'hfd008a8bd86a31ee,64'h91a2d38ed7fe101b,64'he074e519fa557e43,
64'h1efcc283c6a5affb,64'h82949c9da74851ce,64'h9f0e056fd7efb2b8,64'h097467cd50f69617,
64'h8e1170964436ab99,64'h1328b3db16dae060,64'h06de5337752121d1,64'h187bc338b79e92d5,
64'h620ca7689e3b4392,64'h66c109cca2b5225f,64'hd75d0c45ecf13986,64'hfff0000f00100001,
64'h8edb7d6f324d0e5d,64'hbab9048c50810d65,64'hdd4cf314895bf1f8,64'h7546ef77e6fa2fd6,
64'h4394b0dcc558fbf8,64'h544fe11dab2851eb,64'hfe77735095cdcc5c,64'h527757f0fc17202e,
64'h3fb2a0ab3ee3c459,64'hff6cb8b038fddb3b,64'hd34ba3075f23abbd,64'hcb8575222184dc18,
64'ha48693654cee2413,64'hd031d0d956752acf,64'h54ea6dc55923223f,64'hfffffffeffffc001,
64'hba9a67c9f6061e97,64'he8045465c3518f69,64'h8d169c7abff080d4,64'h03a728d6d2abf211,
64'hf7e6141e352d7fd8,64'h14a4e4f13a428e6c,64'hf8702b82bf7d95bc,64'h4ba33e6a87b4b0b8,
64'h708b84b621b55cc4,64'h99459ed8b6d70300,64'h36f299bba9090e88,64'hc3de19c5bcf496a8,
64'h10653b47f1da1c8d,64'h36084e6815a912f5,64'hbae862356789cc2a,64'hff80007f00800001,
64'h76dbeb7d926872e4,64'hd5c8246784086b23,64'hea6798aa4adf8fba,64'haa377bc237d17ead,
64'h1ca586e82ac7dfbe,64'ha27f08ef59428f56,64'hf3bb9a8bae6e62d9,64'h93babf89e0b9016e,
64'hfd95055af71e22c7,64'hfb65c588c7eed9d1,64'h9a5d1840f91d5de2,64'h5c2ba9170c26e0ba,
64'h24349b2f67712093,64'h818e86d0b3a95672,64'ha7536e2cc91911f6,64'hfffffffefffe0001,
64'hd4d33e54b030f4b3,64'h4022a3351a8c7b41,64'h68b4e3d9ff84069c,64'h1d3946b6955f9088,
64'hbf30a0f8a96bfeb9,64'ha5272789d2147360,64'hc3815c1cfbecadd9,64'h5d19f3563da585be,
64'h845c25b40daae61d,64'hca2cf6c9b6b817fc,64'hb794cdde4848743f,64'h1ef0ce33e7a4b53a,
64'h8329da3f8ed0e468,64'hb0427341ad4897a7,64'hd74311b03c4e614b,64'hfc0003ff04000001,
64'hb6df5bef9343971d,64'hae41234220435912,64'h533cc55956fc7dc9,64'h51bbde16be8bf563,
64'he52c3741563efdf0,64'h13f8477fca147aab,64'h9ddcd464737316c1,64'h9dd5fc5305c80b6c,
64'heca82adeb8f11631,64'hdb2e2c4d3f76ce81,64'hd2e8c20bc8eaef0c,64'he15d48ba613705ce,
64'h21a4d97c3b890497,64'h0c7436899d4ab38c,64'h3a9b716b48c88fab,64'hfffffffefff00001,
64'ha699f2ab8187a592,64'h011519aad463da06,64'h45a71ed2fc2034dd,64'he9ca35b4aafc8440,
64'hf98507ca4b5ff5c3,64'h29393c5390a39afb,64'h1c0ae0eddf656ec2,64'he8cf9ab3ed2c2dee,
64'h22e12da46d5730e4,64'h5167b653b5c0bfda,64'hbca66ef74243a1f3,64'hf786719f3d25a9d0,
64'h194ed2007687233c,64'h82139a126a44bd33,64'hba188d87e2730a52,64'he0001fff20000001,
64'hb6fadf819a1cb8e3,64'h72091a16021ac88b,64'h99e62accb7e3ee46,64'h8ddef0b7f45fab16,
64'h2961ba11b1f7ef79,64'h9fc23bfe50a3d558,64'heee6a3279b98b604,64'heeafe29c2e405b5c,
64'h654156fcc788b181,64'hd971626ffbb67402,64'h974610644757785a,64'h0aea45da09b82e69,
64'h0d26cbe2dc4824b7,64'h63a1b44cea559c60,64'hd4db8b5b46447d57,64'hfffffffeff800001,
64'h34cf95610c3d2c8b,64'h08a8cd56a31ed030,64'h2d38f699e101a6e6,64'h4e51adac57e421f9,
64'hcc283e595affae11,64'h49c9e29d851cd7d7,64'he057076efb2b7610,64'h467cd5a669616f69,
64'h17096d246ab9871f,64'h8b3db29fae05fece,64'he53377bf121d0f93,64'hbc338d00e92d4e79,
64'hca769003b43919e0,64'h109cd0975225e994,64'hd0c46c441398528b,64'h0001000000000001,
64'hb7d6fc11d0e5c713,64'h9048d0b310d64455,64'hcf315669bf1f722c,64'h6ef785c3a2fd58ac,
64'h4b0dd08e8fbf7bc7,64'hfe11dff6851eaabc,64'h77351943dcc5b019,64'h757f14e87202dad9,
64'h2a0ab7e93c458c05,64'hcb8b1385ddb3a00a,64'hba3083263abbc2cc,64'h57522ed04dc17348,
64'h69365f16e24125b8,64'h1d0da26a52ace2fd,64'ha6dc5ae03223eab2,64'hfffffffefc000001,
64'ha67cab0961e96457,64'h45466ab518f68180,64'h69c7b4d0080d372f,64'h728d6d64bf210fc6,
64'h6141f2d0d7fd7082,64'h4e4f14ee28e6beb6,64'h02b83b7ed95bb079,64'h33e6ad354b0b7b46,
64'hb84b692355cc38f8,64'h59ed9501702ff66c,64'h299bbdff90e87c91,64'he19c680c496a73c3,
64'h53b48023a1c8cefa,64'h84e684ba912f4ca0,64'h862362269cc29452,64'h0008000000000008,
64'hbeb7e093872e3893,64'h8246859c86b222a4,64'h798ab353f8fb915a,64'h77bc2e2017eac55d,
64'h586e84767dfbde36,64'hf08effbb28f555d9,64'hb9a8ca21e62d80c5,64'habf8a7469016d6c5,
64'h5055bf4ae22c6027,64'h5c589c34ed9d004a,64'hd1841936d5de165b,64'hba9176846e0b9a3e,
64'h49b2f8ba12092dbd,64'he86d1352956717e8,64'h36e2d706911f558b,64'hfffffffee0000001,
64'h33e558500f4b22b3,64'h2a3355aac7b40bfe,64'h4e3da6834069b975,64'h946b6b28f9087e2d,
64'h0a0f9689bfeb840d,64'h7278a7734735f5ae,64'h15c1dbf6cadd83c8,64'h9f3569ab585bda2f,
64'hc25b491fae61c7bb,64'hcf6ca80d817fb35e,64'h4cddeffd8743e487,64'h0ce340694b539e11,
64'h9da4011f0e4677ce,64'h273425d8897a64fc,64'h311b1138e614a28c,64'h0040000000000040,
64'hf5bf04a13971c493,64'h12342ce83591151c,64'hcc559aa2c7dc8acd,64'hbde17103bf562ae5,
64'hc37423b5efdef1ae,64'h8477fde047aaaec1,64'hcd465114316c0623,64'h5fc53a3980b6b623,
64'h82adfa5911630136,64'he2c4e1a96ce8024e,64'h8c20c9bcaef0b2d2,64'hd48bb428705cd1eb,
64'h4d97c5d290496de6,64'h43689a9bab38bf39,64'hb716b83588faac57,64'hfffffffe00000001,
64'h9f2ac2817a591597,64'h519aad573da05fef,64'h71ed341c034dcba6,64'ha35b594bc843f164,
64'h507cb44dff5c2068,64'h93c53b9d39afad6d,64'hae0edfb656ec1e40,64'hf9ab4d5ec2ded174,
64'h12da4903730e3dd2,64'h7b6540720bfd9aea,64'h66ef7fee3a1f2436,64'h671a034a5a9cf088,
64'hed2008fc7233be6c,64'h39a12ec54bd327df,64'h88d889c830a5145f,64'h0200000000000200,
64'hadf82510cb8e2491,64'h91a16741ac88a8e0,64'h62acd51c3ee45662,64'hef0b8822fab15723,
64'h1ba11db57ef78d6a,64'h23bfef063d557604,64'h6a3288a78b603112,64'hfe29d1ce05b5b116,
64'h156fd2cc8b1809ac,64'h16270d5267401269,64'h61064de97785968c,64'ha45da14982e68f52,
64'h6cbe2e96824b6f2e,64'h1b44d4df59c5f9c6,64'hb8b5c1b147d562b3,64'hfffffff700000001,
64'hf956140fd2c8acb4,64'h8cd56abbed02ff76,64'h8f69a0e31a6e5d2d,64'h1adaca63421f8b1b,
64'h83e5a271fae1033e,64'h9e29dcedcd7d6b64,64'h7076fdb7b760f1fb,64'hcd5a6afd16f68b99,
64'h96d2481b9871ee90,64'hdb2a03935fecd74d,64'h377bff74d0f921ad,64'h38d01a55d4e7843d,
64'h690047ea919df359,64'hcd09762b5e993ef7,64'h46c44e458528a2f4,64'h1000000000001000,
64'h6fc1288b5c712483,64'h8d0b3a11644546fc,64'h1566a8e4f722b30d,64'h785c411ed58ab911,
64'hdd08edabf7bc6b50,64'h1dff7832eaabb01f,64'h5194453f5b01888d,64'hf14e8e772dad88a9,
64'hab7e966458c04d60,64'hb1386a933a009348,64'h08326f4ebc2cb45d,64'h22ed0a5117347a8b,
64'h65f174b7125b796d,64'hda26a6face2fce30,64'hc5ae0d8f3eab1593,64'hffffffbf00000001,
64'hcab0a08596456599,64'h66ab55e36817fbac,64'h7b4d071cd372e964,64'hd6d6531a10fc58d8,
64'h1f2d1393d70819ec,64'hf14ee7726beb5b1c,64'h83b7edc0bb078fd5,64'h6ad357eeb7b45cc2,
64'hb69240e0c38f747c,64'hd9501ca0ff66ba62,64'hbbdffba787c90d67,64'hc680d2afa73c21e7,
64'h48023f578cef9ac5,64'h684bb160f4c9f7b2,64'h3622722e2945179e,64'h8000000000008000,
64'h7e09445de3892415,64'h6859d08f222a37dc,64'hab354727b9159868,64'hc2e208f9ac55c885,
64'he8476d65bde35a7a,64'heffbc197555d80f8,64'h8ca229fcd80c4466,64'h8a7473c06d6c4541,
64'h5bf4b327c6026afb,64'h89c3549ed0049a3b,64'h41937a75e165a2e8,64'h17685289b9a3d457,
64'h2f8ba5bb92dbcb65,64'hd13537dc717e717a,64'h2d706c7ff558ac92,64'hfffffdff00000001,
64'h55850432b22b2cc2,64'h355aaf1e40bfdd5d,64'hda6838e99b974b1d,64'hb6b298d687e2c6ba,
64'hf9689c9eb840cf60,64'h8a773b9a5f5ad8d9,64'h1dbf6e09d83c7ea4,64'h569abf78bda2e60d,
64'hb492070b1c7ba3db,64'hca80e50dfb35d30a,64'hdeffdd413e486b33,64'h3406958339e10f32,
64'h4011fabe677cd626,64'h425d8b0aa64fbd8d,64'hb11391724a28bcef,64'h000000040003fffc,
64'hf04a22f21c4920a5,64'h42ce847c1151bedd,64'h59aa3942c8acc33b,64'h171047d362ae4422,
64'h423b6b34ef1ad3c9,64'h7fde0cc1aaec07b9,64'h65114feac062232c,64'h53a39e076b622a04,
64'hdfa59940301357d6,64'h4e1aa4fa8024d1d4,64'h0c9bd3b10b2d173e,64'hbb42944dcd1ea2b8,
64'h7c5d2ddd96de5b27,64'h89a9bee98bf38bca,64'h6b836400aac5648f,64'hffffefff00000001,
64'hac2821979159660e,64'haad578f305feeae7,64'hd341c752dcba58e2,64'hb594c6b93f1635cb,
64'hcb44e4fcc2067af9,64'h53b9dcd6fad6c6c4,64'hedfb704ec1e3f520,64'hb4d5fbc7ed173066,
64'ha490385de3dd1ed3,64'h54072875d9ae984a,64'hf7feea0ff2435992,64'ha034ac1acf08798f,
64'h008fd5f53be6b12e,64'h12ec5857327dec66,64'h889c8b975145e773,64'h00000020001fffe0,
64'h82511797e2490521,64'h167423e28a8df6e6,64'hcd51ca18456619d6,64'hb8823e9b15722110,
64'h11db59a978d69e46,64'hfef0661057603dc5,64'h288a7f590311195d,64'h9d1cf03d5b11501e,
64'hfd2cca07809abeaa,64'h70d527d601268e9e,64'h64de9d885968b9f0,64'hda14a27368f515bb,
64'he2e96eefb6f2d935,64'h4d4df7505f9c5e4c,64'h5c1b2008562b2475,64'hffff7fff00000001,
64'h61410cc18acb306b,64'h56abc79d2ff75733,64'h9a0e3a9ce5d2c70a,64'haca635cef8b1ae53,
64'h5a2727ec1033d7c2,64'h9dcee6b9d6b6361e,64'h6fdb827d0f1fa8f9,64'ha6afde4468b9832b,
64'h2481c2f41ee8f693,64'ha03943b0cd74c24e,64'hbff75086921acc89,64'h01a560db7843cc73,
64'h047eafa9df358970,64'h9762c2b993ef6330,64'h44e45cbe8a2f3b94,64'h0000010000ffff00,
64'h1288bcc312482904,64'hb3a11f14546fb730,64'h6a8e50c82b30ceaa,64'hc411f4ddab91087b,
64'h8edacd4bc6b4f230,64'hf7833089bb01ee21,64'h4453fac91888cae7,64'he8e781eed88a80ec,
64'he966504304d5f549,64'h86a93eb3093474ed,64'h26f4ec45cb45cf7d,64'hd0a513a147a8add2,
64'h174b7784b796c9a1,64'h6a6fba84fce2f25e,64'he0d90044b15923a6,64'hfffbffff00000001,
64'h0a08660f56598355,64'hb55e3ceb7fbab996,64'hd071d4eb2e96384c,64'h6531ae7cc58d7293,
64'hd1393f62819ebe0e,64'hee7735d2b5b1b0ec,64'h7edc13eb78fd47c5,64'h357ef22845cc1953,
64'h240e17a1f747b497,64'h01ca1d8b6ba6126b,64'hffba843990d66443,64'h0d2b06dbc21e6398,
64'h23f57d4ef9ac4b80,64'hbb1615d09f7b197c,64'h2722e5f65179dc9e,64'h0000080007fff800,
64'h9445e61892414820,64'h9d08f8a7a37db97b,64'h547286445986754d,64'h208fa6f35c8843d2,
64'h76d66a6235a7917c,64'hbc198454d80f7101,64'h229fd64ac4465736,64'h473c0f7dc4540759,
64'h4b32821f26afaa41,64'h3549f59c49a3a764,64'h37a7622f5a2e7be7,64'h85289d103d456e8a,
64'hba5bbc25bcb64d08,64'h537dd42ae71792ed,64'h06c8022c8ac91d29,64'hffdfffff00000001,
64'h5043307ab2cc1aa8,64'haaf1e760fdd5ccab,64'h838ea75f74b1c25a,64'h298d73e92c6b9495,
64'h89c9fb1a0cf5f06a,64'h73b9ae9cad8d8759,64'hf6e09f5ec7ea3e25,64'habf791432e60ca97,
64'h2070bd10ba3da4b7,64'h0e50ec5b5d309358,64'hfdd421d386b32211,64'h695836de10f31cc0,
64'h1fabea78cd625bff,64'hd8b0ae89fbd8cbdb,64'h39172fb38bcee4ef,64'h000040003fffc000,
64'ha22f30c8920a40fc,64'he847c5411bedcbd4,64'ha3943224cc33aa66,64'h047d379be4421e8f,
64'hb6b35314ad3c8bdd,64'he0cc22abc07b8803,64'h14feb2572232b9af,64'h39e07bf022a03ac6,
64'h599410fb357d5206,64'haa4face34d1d3b1f,64'hbd3b117bd173df37,64'h2944e885ea2b744c,
64'hd2dde132e5b2683b,64'h9beea15938bc9766,64'h364011645648e948,64'hfeffffff00000001,
64'h821983d79660d53e,64'h578f3b0ceeae6553,64'h1c753affa58e12cc,64'h4c6b9f4a635ca4a7,
64'h4e4fd8d467af834c,64'h9dcd74e86c6c3ac5,64'hb704fafd3f51f121,64'h5fbc8a1e730654b3,
64'h0385e886d1ed25b7,64'h728762dae9849ac0,64'heea10ea335991081,64'h4ac1b6f38798e5fd,
64'hfd5f53c66b12dff8,64'hc5857455dec65ed2,64'hc8b97d9d5e772777,64'h00020001fffe0000,
64'h11798649905207db,64'h423e2a0fdf6e5e99,64'h1ca1912b619d532b,64'h23e9bcdf2210f478,
64'hb59a98aa69e45ee3,64'h0661156503dc4011,64'ha7f592b91195cd78,64'hcf03df821501d62f,
64'hcca087dbabea902e,64'h527d671f68e9d8f3,64'he9d88be38b9ef9b3,64'h4a274430515ba25f,
64'h96ef099d2d9341d2,64'hdf750acdc5e4bb2c,64'hb2008b23b2474a3f,64'hf7ffffff00000001,
64'h10cc1ec0b306a9ec,64'hbc79d86975732a96,64'he3a9d7fd2c709660,64'h635cfa551ae52536,
64'h727ec6a53d7c1a5e,64'hee6ba7476361d624,64'hb827d7eefa8f8903,64'hfde450f59832a596,
64'h1c2f44368f692db8,64'h943b16da4c24d5fd,64'h75087520acc88401,64'h560db79e3cc72fe6,
64'heafa9e3a5896ffb9,64'h2c2ba2b4f632f68a,64'h45cbecf0f3b93bb2,64'h0010000ffff00000,
64'h8bcc324c82903ed8,64'h11f15080fb72f4c6,64'he50c895b0cea9958,64'h1f4de6fa1087a3bf,
64'hacd4c5584f22f713,64'h3308ab281ee20088,64'h3fac95cd8cae6bbb,64'h781efc16a80eb172,
64'h65043ee35f54816a,64'h93eb38fd474ec796,64'h4ec45f235cf7cd91,64'h513a21848add12f6,
64'hb7784ced6c9a0e8c,64'hfba856742f25d95a,64'h90045922923a51f3,64'hbfffffff00000001,
64'h8660f60598354f60,64'he3cec350ab9954ab,64'h1d4ebff06384b2f9,64'h1ae7d2abd72929ad,
64'h93f6352cebe0d2ed,64'h735d3a421b0eb119,64'hc13ebf7cd47c4813,64'hef2287b3c1952ca9,
64'he17a21b47b496dc0,64'ha1d8b6d66126afe4,64'ha843a90866442005,64'hb06dbcf3e6397f2e,
64'h57d4f1d9c4b7fdc1,64'h615d15a8b197b44f,64'h2e5f67899dc9dd8e,64'h0080007fff800000,
64'h5e6192681481f6bc,64'h8f8a8407db97a630,64'h28644adf6754cab9,64'hfa6f37d0843d1df8,
64'h66a62ac77917b893,64'h98455941f710043f,64'hfd64ae6d65735dd7,64'hc0f7e0b840758b8d,
64'h2821f71dfaa40b4d,64'h9f59c7ee3a763cac,64'h7622f91ce7be6c86,64'h89d10c2656e897ae,
64'hbbc2677064d0745b,64'hdd42b3a8792ecac9,64'h8022c91891d28f94,64'hfffffffd00000003,
64'h3307b030c1aa7afc,64'h1e761a8c5ccaa551,64'hea75ff831c2597c8,64'hd73e955eb9494d68,
64'h9fb1a96b5f069764,64'h9ae9d213d87588c5,64'h09f5fbeca3e24092,64'h79143da50ca96541,
64'h0bd10daada4b6df9,64'h0ec5b6b809357f1b,64'h421d484832210023,64'h836de7a431cbf96b,
64'hbea78ed025bfee06,64'h0ae8ad488cbda275,64'h72fb3c4dee4eec6f,64'h040003fffc000000,
64'hf30c9342a40fb5de,64'h7c542042dcbd317c,64'h432256fc3aa655c7,64'hd379be8b21e8efb9,
64'h3531563ec8bdc495,64'hc22aca13b88021f4,64'heb2573722b9aeeb1,64'h07bf05c803ac5c62,
64'h410fb8f0d5205a67,64'hface3f75d3b1e55c,64'hb117c8ea3df3642d,64'h4e886136b744bd6c,
64'hde133b882683a2d3,64'hea159d49c9765642,64'h011648c88e947c9c,64'hffffffef00000011,
64'h983d81870d53d7df,64'hf3b0d462e6552a88,64'h53affc1fe12cbe39,64'hb9f4aafbca4a6b3a,
64'hfd8d4b5ef834bb1c,64'hd74e90a2c3ac4624,64'h4fafdf651f120490,64'hc8a1ed2b654b2a05,
64'h5e886d56d25b6fc8,64'h762db5c049abf8d8,64'h10ea424391080116,64'h1b6f3d258e5fcb54,
64'hf53c76862dff702b,64'h57456a4465ed13a8,64'h97d9e27272776375,64'h20001fffe0000000,
64'h98649a1c207daee9,64'he2a10219e5e98bdd,64'h1912b7e3d532ae36,64'h9bcdf45f0f477dc2,
64'ha98ab1f745ee24a7,64'h115650a3c4010f9a,64'h592b9b985cd77581,64'h3df82e401d62e310,
64'h087dc788a902d336,64'hd671fbb59d8f2ad9,64'h88be4756ef9b2163,64'h744309b7ba25eb5e,
64'hf099dc47341d1692,64'h50acea554bb2b209,64'h08b2464474a3e4e0,64'hffffff7f00000081,
64'hc1ec0c3c6a9ebef4,64'h9d86a31e32a95439,64'h9d7fe1010965f1c6,64'hcfa557e3525359cb,
64'hec6a5afec1a5d8d9,64'hba74851c1d62311a,64'h7d7efb2af890247e,64'h450f69612a595022,
64'hf4436ab892db7e3e,64'hb16dae054d5fc6bd,64'h8752121c884008b0,64'hdb79e92c72fe5aa0,
64'ha9e3b4386ffb8151,64'hba2b52252f689d3e,64'hbecf139793bb1ba4,64'h0000ffffffffffff,
64'hc324d0e503ed7744,64'h150810d62f4c5ee1,64'hc895bf1ea99571b0,64'hde6fa2fc7a3bee0c,
64'h4c558fbf2f712533,64'h8ab2851e20087cd0,64'hc95cdcc4e6bbac06,64'hefc17201eb17187f,
64'h43ee3c45481699b0,64'hb38fddb2ec7956c2,64'h45f23abb7cd90b14,64'ha2184dc0d12f5aed,
64'h84cee240a0e8b489,64'h856752ac5d959046,64'h45923223a51f2700,64'hfffffbff00000401,
64'h0f6061e954f5f79a,64'hec3518f5954aa1c4,64'hebff080c4b2f8e2c,64'h7d2abf20929ace52,
64'h6352d7fd0d2ec6c1,64'hd3a428e5eb1188cb,64'hebf7d95ac48123ed,64'h287b4b0b52ca810e,
64'ha21b55cb96dbf1e9,64'h8b6d702f6afe35e3,64'h3a9090e84200457c,64'hdbcf496997f2d4fa,
64'h4f1da1c87fdc0a83,64'hd15a912e7b44e9eb,64'hf6789cc19dd8dd1b,64'h0007fffffffffff8,
64'h1926872e1f6bba1a,64'ha84086b17a62f708,64'h44adf8fb4cab8d7a,64'hf37d17e9d1df705a,
64'h62ac7dfb7b892996,64'h559428f50043e67c,64'h4ae6e62d35dd602a,64'h7e0b901658b8c3f1,
64'h1f71e22c40b4cd7e,64'h9c7eed9c63cab60b,64'h2f91d5dde6c8589e,64'h10c26e0b897ad763,
64'h267712090745a444,64'h2b3a9566ecac822c,64'h2c91911f28f937fe,64'hffffdfff00002001,
64'h7b030f4aa7afbcd0,64'h61a8c7b3aa550e19,64'h5ff84069597c7159,64'he955f90794d6728d,
64'h1a96bfeb69763605,64'h9d214735588c4652,64'h5fbecadd24091f61,64'h43da585b9654086f,
64'h10daae61b6df8f43,64'h5b6b817f57f1af14,64'hd484874310022bdf,64'hde7a4b52bf96a7ca,
64'h78ed0e45fee05416,64'h8ad48979da274f52,64'hb3c4e613eec6e8d1,64'h003fffffffffffc0,
64'hc9343970fb5dd0d0,64'h42043590d317b83b,64'h256fc7dc655c6bce,64'h9be8bf558efb82c9,
64'h1563efdedc494cad,64'haca147aa021f33de,64'h5737316baeeb014e,64'hf05c80b5c5c61f85,
64'hfb8f116205a66bf0,64'he3f76ce71e55b054,64'h7c8eaef03642c4ef,64'h8613705c4bd6bb18,
64'h33b890493a2d221f,64'h59d4ab386564115f,64'h648c88fa47c9bfef,64'hfffeffff00010001,
64'hd8187a583d7de67d,64'h0d463da052a870c5,64'hffc2034ccbe38ac6,64'h4aafc843a6b39461,
64'hd4b5ff5b4bb1b028,64'he90a39aec462328c,64'hfdf656eb2048fb06,64'h1ed2c2deb2a04376,
64'h86d5730db6fc7a18,64'hdb5c0bfcbf8d789e,64'ha4243a1e80115ef2,64'hf3d25a9bfcb53e4a,
64'hc7687232f702a0ad,64'h56a44bd2d13a7a8c,64'h9e2730a476374683,64'h01fffffffffffe00,
64'h49a1cb8ddaee867a,64'h1021ac8898bdc1d6,64'h2b7e3ee42ae35e6f,64'hdf45fab077dc1644,
64'hab1f7ef6e24a6568,64'h650a3d5510f99eeb,64'hb9b98b5f77580a6e,64'h82e405b52e30fc21,
64'hdc788b172d335f79,64'h1fbb673ff2ad8299,64'he4757784b2162775,64'h309b82e65eb5d8bc,
64'h9dc4824ad16910f7,64'hcea559c52b208af6,64'h246447d53e4dff75,64'hfff7ffff00080001,
64'hc0c3d2c7ebef33e2,64'h6a31ed0295438628,64'hfe101a6d5f1c5629,64'h557e421f359ca306,
64'ha5affae05d8d813a,64'h4851cd7d23119459,64'hefb2b7600247d829,64'hf69616f595021bb0,
64'h36ab9871b7e3d0bc,64'hdae05febfc6bc4ea,64'h2121d0f9008af78b,64'h9e92d4e6e5a9f249,
64'h3b43919db8150562,64'hb5225e9889d3d45e,64'hf1398527b1ba3414,64'h0ffffffffffff000,
64'h4d0e5c70d77433ce,64'h810d6444c5ee0eb0,64'h5bf1f722571af377,64'hfa2fd589bee0b21a,
64'h58fbf7bc12532b3b,64'h2851eaab87ccf755,64'hcdcc5b00bac0536b,64'h17202dad7187e104,
64'he3c458bf699afbc2,64'hfddb39ff956c14c8,64'h23abbc2c90b13ba1,64'h84dc1733f5aec5df,
64'hee24125a8b4887b4,64'h752ace2f590457aa,64'h23223eaaf26ffba7,64'hffbfffff00400001
};
  //------------------------
  // 512
  //------------------------
  localparam [2*512-1:0][63:0] NTT_GF64_BWD_WDIV_N512_PHI_L = {
64'ha31ed02f5438627a,64'h57e421f859ca305b,64'h851cd7d63119458c,64'h69616f685021baf1,
64'hae05feccc6bc4e93,64'he92d4e775a9f2487,64'h5225e9939d3d45d5,64'h00000000fffeffff,
64'h10d644545ee0eaf8,64'ha2fd58aaee0b2191,64'h851eaaba7ccf754e,64'h7202dad8187e103f,
64'hddb3a00856c14c71,64'h4dc173475aec5de8,64'h52ace2fc90457a99,64'hfbffffff04000001,
64'h18f6817fa1c313cb,64'hbf210fc4ce5182d6,64'h28e6beb588ca2c5c,64'h4b0b7b45810dd785,
64'h702ff66b35e27493,64'h496a73c1d4f92431,64'h912f4c9ee9ea2ea6,64'h00000007fff7fff8,
64'h86b222a2f70757c0,64'h17eac55c70590c83,64'h28f555d7e67baa6c,64'h9016d6c3c3f081f5,
64'hed9d0048b60a6382,64'h6e0b9a3cd762ef3e,64'h956717e6822bd4c6,64'hdfffffff20000001,
64'hc7b40bfd0e189e58,64'hf9087e2b728c16ab,64'h4735f5ad465162df,64'h585bda2e086ebc26,
64'h817fb35caf13a495,64'h4b539e10a7c92186,64'h897a64fb4f51752c,64'h0000003fffbfffc0,
64'h3591151bb83abdfc,64'hbf562ae382c86418,64'h47aaaec033dd535f,64'h80b6b6221f840fa4,
64'h6ce8024cb0531c09,64'h705cd1e9bb1779ed,64'hab38bf38115ea62c,64'h0000000000000001,
64'h3da05fee70c4f2ba,64'hc843f1629460b551,64'h39afad6c328b16f6,64'hc2ded1724375e12e,
64'h0bfd9ae9789d24a4,64'h5a9cf0873e490c2e,64'h4bd327de7a8ba95c,64'h000001fffdfffe00,
64'hac88a8dec1d5efdf,64'hfab15721164320bb,64'h3d5576039eea9af6,64'h05b5b114fc207d1c,
64'h674012688298e045,64'h82e68f50d8bbcf65,64'h59c5f9c58af5315b,64'h0000000000000008,
64'hed02ff74862795cf,64'h421f8b1aa305aa82,64'hcd7d6b629458b7af,64'h16f68b981baf096a,
64'h5fecd74bc4e92520,64'hd4e7843bf248616e,64'h5e993ef5d45d4ade,64'h00000fffeffff000,
64'h644546fb0eaf7ef3,64'hd58ab90fb21905d1,64'heaabb01df754d7af,64'h2dad88a7e103e8e0,
64'h3a00934714c70225,64'h17347a8ac5de7b24,64'hce2fce2e57a98ad6,64'h0000000000000040,
64'h6817fbab313cae71,64'h10fc58d7182d540e,64'h6beb5b1aa2c5bd72,64'hb7b45cc0dd784b50,
64'hff66ba60274928fe,64'ha73c21e592430b6a,64'hf4c9f7b0a2ea56ee,64'h00007fff7fff8000,
64'h222a37db757bf795,64'hac55c88390c82e82,64'h555d80f6baa6bd71,64'h6d6c4540081f46ff,
64'hd0049a39a6381127,64'hb9a3d4562ef3d920,64'h717e7178bd4c56aa,64'h0000000000000200,
64'h40bfdd5c89e57385,64'h87e2c6b8c16aa070,64'h5f5ad8d8162deb8d,64'hbda2e60bebc25a7b,
64'hfb35d3083a4947e9,64'h39e10f3192185b4b,64'ha64fbd8c1752b769,64'h0003fffbfffc0000,
64'h1151bedcabdfbca7,64'h62ae44218641740b,64'haaec07b7d535eb86,64'h6b622a0340fa37f5,
64'h8024d1d331c08932,64'hcd1ea2b6779ec8fb,64'h8bf38bc8ea62b54d,64'h0000000000001000,
64'h05feeae64f2b9c26,64'h3f1635ca0b55037c,64'hfad6c6c2b16f5c66,64'hed1730645e12d3d3,
64'hd9ae9848d24a3f41,64'hcf08798d90c2da57,64'h327dec65ba95bb43,64'h001fffdfffe00000,
64'h8a8df6e55efde538,64'h1572210f320ba055,64'h57603dc3a9af5c2b,64'h5b11501d07d1bfa5,
64'h01268e9d8e04498c,64'h68f515b9bcf647d2,64'h5f9c5e4b5315aa64,64'h0000000000008000,
64'h2ff75732795ce130,64'hf8b1ae515aa81bdf,64'hd6b6361c8b7ae329,64'h68b98329f0969e91,
64'hcd74c24c9251fa02,64'h7843cc728616d2b2,64'h93ef632ed4adda17,64'h00fffeffff000000,
64'h546fb72ef7ef29bc,64'hab910879905d02a8,64'hbb01ee1f4d7ae156,64'hd88a80ea3e8dfd26,
64'h093474ec70224c60,64'h47a8add0e7b23e8d,64'hfce2f25c98ad531e,64'h0000000000040000,
64'h7fbab994cae7097f,64'hc58d7291d540def1,64'hb5b1b0ea5bd71942,64'h45cc195284b4f485,
64'h6ba6126a928fd00a,64'hc21e639730b6958d,64'h9f7b197aa56ed0b4,64'h07fff7fff8000000,
64'ha37db979bf794dde,64'h5c8843d182e8153b,64'hd80f70ff6bd70aab,64'hc4540757f46fe92a,
64'h49a3a76381126300,64'h3d456e893d91f466,64'he71792ebc56a98e9,64'h0000000000200000,
64'hfdd5cca957384bf5,64'h2c6b9494aa06f782,64'had8d8757deb8ca0b,64'h2e60ca9625a7a426,
64'h5d309357947e804d,64'h10f31cbf85b4ac62,64'hfbd8cbd92b76859c,64'h3fffbfffc0000000,
64'h1bedcbd2fbca6eeb,64'he4421e8e1740a9d6,64'hc07b88015eb85552,64'h22a03ac5a37f494a,
64'h4d1d3b1e089317fe,64'hea2b744aec8fa32f,64'h38bc97652b54c741,64'h0000000001000000,
64'heeae6551b9c25fa1,64'h635ca4a65037bc0f,64'h6c6c3ac3f5c65053,64'h730654b22d3d212f,
64'he9849abea3f40266,64'h8798e5fc2da56310,64'hdec65ed05bb42cd9,64'hfffdfffeffffffff,
64'hdf6e5e97de537758,64'h2210f477ba054ea9,64'h03dc4010f5c2aa8a,64'h1501d62e1bfa4a4f,
64'h68e9d8f24498bfee,64'h515ba25e647d1971,64'hc5e4bb2a5aa63a07,64'h0000000008000000,
64'h75732a94ce12fd01,64'h1ae5253581bde075,64'h6361d622ae328295,64'h9832a59469e90975,
64'h4c24d5fc1fa01329,64'h3cc72fe56d2b187c,64'hf632f688dda166c2,64'hffeffffefffffff1,
64'hfb72f4c4f29bbaba,64'h1087a3bed02a7547,64'h1ee20087ae155450,64'ha80eb170dfd25278,
64'h474ec79524c5ff6d,64'h8add12f523e8cb86,64'h2f25d958d531d032,64'h0000000040000000,
64'hab9954a97097e805,64'hd72929ac0def03a8,64'h1b0eb118719414a5,64'hc1952ca74f484ba4,
64'h6126afe2fd009946,64'he6397f2c6958c3df,64'hb197b44ded0b3609,64'hff7ffffeffffff81,
64'hdb97a62e94ddd5c9,64'h843d1df68153aa38,64'hf710043d70aaa280,64'h40758b8bfe9293bb,
64'h3a763cab262ffb66,64'h56e897ad1f465c2c,64'h792ecac7a98e818f,64'h0000000200000000,
64'h5ccaa55084bf4023,64'hb9494d666f781d3a,64'hd87588c38ca0a528,64'h0ca965407a425d1a,
64'h09357f1ae804ca2d,64'h31cbf96a4ac61ef1,64'h8cbda2746859b043,64'hfbfffffefffffc01,
64'hdcbd317aa6eeae42,64'h21e8efb80a9d51bc,64'hb88021f2855513f9,64'h03ac5c61f4949dd6,
64'hd3b1e55a317fdb2f,64'hb744bd6afa32e15e,64'hc97656404c740c75,64'h0000001000000000,
64'he6552a8625fa0116,64'hca4a6b387bc0e9cb,64'hc3ac46226505293a,64'h654b2a03d212e8d0,
64'h49abf8d740265168,64'h8e5fcb535630f787,64'h65ed13a742cd8214,64'hdffffffeffffe001,
64'he5e98bdb3775720a,64'h0f477dc154ea8ddf,64'hc4010f992aa89fc3,64'h1d62e30fa4a4eeb0,
64'h9d8f2ad78bfed972,64'hba25eb5cd1970aeb,64'h4bb2b20863a063a2,64'h0000008000000000,
64'h32a954382fd008a9,64'h525359c9de074e52,64'h1d623119282949ca,64'h2a5950219097467d,
64'h4d5fc6bc01328b3e,64'h72fe5a9eb187bc34,64'h2f689d3d166c109d,64'hfffffffdffff0002,
64'h2f4c5ee0bbab9049,64'h7a3bee0aa7546ef8,64'h20087ccf5544fe12,64'heb17187d25277580,
64'hec7956c05ff6cb8c,64'hd12f5aeb8cb85753,64'h5d9590451d031d0e,64'h0000040000000000,
64'h954aa1c27e804547,64'h929ace50f03a728e,64'heb1188c9414a4e50,64'h52ca810d84ba33e7,
64'h6afe35e2099459ee,64'h97f2d4f88c3de19d,64'h7b44e9e9b36084e7,64'hfffffff6fff80009,
64'h7a62f706dd5c8247,64'hd1df70583aa377bd,64'h0043e67baa27f08f,64'h58b8c3f0293babf9,
64'h63cab609ffb65c59,64'h897ad76265c2ba92,64'hecac822ae818e86e,64'h0000200000000000,
64'haa550e17f4022a34,64'h94d6728b81d3946c,64'h588c46510a527279,64'h9654086e25d19f36,
64'h57f1af134ca2cf6d,64'hbf96a7c861ef0ce4,64'hda274f509b042735,64'hffffffbeffc00041,
64'hd317b839eae41235,64'h8efb82c7d51bbde2,64'h021f33dd513f8478,64'hc5c61f8349dd5fc6,
64'h1e55b052fdb2e2c5,64'h4bd6bb172e15d48c,64'h6564115e40c74369,64'h0001000000000000,
64'h52a870c4a011519b,64'ha6b394600e9ca35c,64'hc462328a529393c6,64'hb2a043752e8cf9ac,
64'hbf8d789c65167b66,64'hfcb53e480f78671b,64'hd13a7a8ad82139a2,64'hfffffdfefe000201,
64'h98bdc1d5572091a2,64'h77dc1642a8ddef0c,64'h10f99eea89fc23c0,64'h2e30fc204eeafe2a,
64'hf2ad8297ed971628,64'h5eb5d8bb70aea45e,64'h2b208af5063a1b45,64'h0008000000000000,
64'h95438627008a8cd6,64'h359ca30574e51adb,64'h23119458949c9e2a,64'h95021bae7467cd5b,
64'hfc6bc4e828b3db2b,64'he5a9f2477bc338d1,64'h89d3d45cc109cd0a,64'hffffeffef0001001,
64'hc5ee0eaeb9048d0c,64'hbee0b21846ef785d,64'h87ccf7544fe11e00,64'h7187e1037757f14f,
64'h956c14c66cb8b139,64'hf5aec5dd857522ee,64'h590457a931d0da27,64'h0040000000000000,
64'haa1c313c045466ac,64'hace5182ca728d6d7,64'h188ca2c5a4e4f14f,64'ha810dd77a33e6ad4,
64'he35e2748459ed951,64'h2d4f9242de19c681,64'h4e9ea2ea084e684c,64'hffff7ffe80008001,
64'h2f70757bc824685a,64'hf70590c7377bc2e3,64'h3e67baa67f08effc,64'h8c3f081ebabf8a75,
64'hab60a63765c589c4,64'had762ef32ba91769,64'hc822bd4b8e86d136,64'h0200000000000000,
64'h50e189e522a3355b,64'h6728c16a3946b6b3,64'hc465162d27278a78,64'h4086ebc219f3569b,
64'h1af13a492cf6ca81,64'h6a7c9217f0ce3407,64'h74f517524273425e,64'hfffbfffb00040001,
64'h7b83abdf412342cf,64'hb82c8640bbde1711,64'hf33dd534f8477fdf,64'h61f840f9d5fc53a4,
64'h5b0531c02e2c4e1b,64'h6bb1779e5d48bb43,64'h4115ea62743689aa,64'h1000000000000000,
64'h870c4f2b1519aad6,64'h39460b54ca35b595,64'h2328b16f393c53ba,64'h04375e12cf9ab4d6,
64'hd789d24967b65408,64'h53e490c28671a035,64'ha7a8ba95139a12ed,64'hffdfffdf00200001,
64'hdc1d5efd091a1675,64'hc164320adef0b883,64'h99eea9aec23bfef1,64'h0fc207d1afe29d1d,
64'hd8298e03716270d6,64'h5d8bbcf5ea45da15,64'h08af5315a1b44d4e,64'h8000000000000000,
64'h3862795ca8cd56ac,64'hca305aa751adaca7,64'h19458b7ac9e29dcf,64'h21baf0967cd5a6b0,
64'hbc4e92513db2a03a,64'h9f248616338d01a6,64'h3d45d4ad9cd09763,64'hfefffeff01000001,
64'he0eaf7ee48d0b3a2,64'h0b21905cf785c412,64'hcf754d7a11dff784,64'h7e103e8d7f14e8e8,
64'hc14c70218b1386aa,64'hec5de7b1522ed0a6,64'h457a98ad0da26a70,64'h00000003fffffffc,
64'hc313cae6466ab55f,64'h5182d5408d6d6532,64'hca2c5bd64f14ee78,64'h0dd784b4e6ad357f,
64'he274928eed9501cb,64'hf92430b59c680d2c,64'hea2ea56de684bb17,64'hf7fff7ff08000001,
64'h0757bf7946859d09,64'h590c82e7bc2e2090,64'h7baa6bd68effbc1a,64'hf081f46ef8a7473d,
64'h0a638112589c354a,64'h62ef3d9191768529,64'h2bd4c56a6d13537e,64'h0000001fffffffe0,
64'h189e57383355aaf2,64'h8c16aa066b6b298e,64'h5162deb878a773ba,64'h6ebc25a73569abf8,
64'h13a4947e6ca80e51,64'hc92185b3e3406959,64'h51752b763425d8b1,64'hbfffbfff40000001,
64'h3abdfbca342ce848,64'hc864173fe171047e,64'hdd535eb777fde0cd,64'h840fa37ec53a39e1,
64'h531c0892c4e1aa50,64'h1779ec8f8bb42945,64'h5ea62b54689a9bef,64'h000000ffffffff00,
64'hc4f2b9c19aad5790,64'h60b550375b594c6c,64'h8b16f5c5c53b9dce,64'h75e12d3cab4d5fbd,
64'h9d24a3f365407288,64'h490c2da51a034ac2,64'h8ba95bb3a12ec586,64'hfffdffff00000003,
64'hd5efde52a167423f,64'h4320ba050b8823ea,64'hea9af5c1bfef0662,64'h207d1bfa29d1cf04,
64'h98e04498270d527e,64'hbbcf647c5da14a28,64'hf5315aa544d4df76,64'h000007fffffff800,
64'h2795ce12d56abc7a,64'h05aa81bddaca635d,64'h58b7ae3229dcee6c,64'haf0969e85a6afde5,
64'he9251f9f2a03943c,64'h48616d2ad01a560e,64'h5d4adda109762c2c,64'hffefffff00000011,
64'haf7ef29b0b3a11f2,64'h1905d02a5c411f4e,64'h54d7ae14ff783309,64'h03e8dfd24e8e781f,
64'hc70224c5386a93ec,64'hde7b23e7ed0a513b,64'ha98ad53126a6fba9,64'h00003fffffffc000,
64'h3cae7097ab55e3cf,64'h2d540deed6531ae8,64'hc5bd71934ee7735e,64'h784b4f47d357ef23,
64'h4928fd00501ca1d9,64'h430b695880d2b06e,64'hea56ed0a4bb1615e,64'hff7fffff00000081,
64'h7bf794dd59d08f8b,64'hc82e8152e208fa70,64'ha6bd70a9fbc19846,64'h1f46fe927473c0f8,
64'h3811262fc3549f5a,64'hf3d91f45685289d2,64'h4c56a98e3537dd43,64'h0001fffffffe0000,
64'he57384be5aaf1e77,64'h6aa06f77b298d73f,64'h2deb8ca0773b9aea,64'hc25a7a419abf7915,
64'h4947e80480e50ec6,64'h185b4ac60695836e,64'h52b768595d8b0ae9,64'hfbffffff00000401,
64'hdfbca6edce847c55,64'h41740a9d1047d37a,64'h35eb8554de0cc22b,64'hfa37f493a39e07c0,
64'hc089317f1aa4facf,64'h9ec8fa3242944e89,64'h62b54c73a9beea16,64'h000ffffffff00000,
64'h2b9c25f9d578f3b1,64'h55037bc094c6b9f5,64'h6f5c6504b9dcd74f,64'h12d3d212d5fbc8a2,
64'h4a3f40260728762e,64'hc2da563034ac1b70,64'h95bb42ccec585746,64'hdfffffff00002001,
64'hfde537747423e2a2,64'h0ba054ea823e9bce,64'haf5c2aa7f0661157,64'hd1bfa4a41cf03df9,
64'h04498bfed527d672,64'hf647d19614a27444,64'h15aa63a04df750ad,64'h007fffffff800000,
64'h5ce12fcfabc79d87,64'ha81bde06a635cfa6,64'h7ae32828cee6ba75,64'h969e9096afde4510,
64'h51fa01323943b16e,64'h16d2b187a560db7a,64'hadda166b62c2ba2c,64'hfffffffe00010002,
64'hef29bbaaa11f1509,64'h5d02a75411f4de70,64'h7ae1554483308ab3,64'h8dfd2526e781efc2,
64'h224c5ff6a93eb390,64'hb23e8cb7a513a219,64'had531d026fba8568,64'h03fffffffc000000,
64'he7097e7f5e3cec36,64'h40def03a31ae7d2b,64'hd71941497735d3a5,64'hb4f484b97ef2287c,
64'h8fd00993ca1d8b6e,64'hb6958c3d2b06dbd0,64'h6ed0b3601615d15b,64'hfffffff700080009,
64'h794ddd5c08f8a841,64'he8153aa28fa6f37e,64'hd70aaa2719845595,64'h6fe9293b3c0f7e0c,
64'h1262ffb649f59c7f,64'h91f465c2289d10c3,64'h6a98e8187dd42b3b,64'h1fffffffe0000000,
64'h384bf401f1e761a9,64'h06f781d38d73e956,64'hb8ca0a51b9ae9d22,64'ha7a425d0f79143db,
64'h7e804ca250ec5b6c,64'hb4ac61ee5836de7b,64'h76859b03b0ae8ad5,64'hffffffbf00400041,
64'hca6eeae347c54205,64'h40a9d51b7d379be9,64'hb855513ecc22aca2,64'h7f4949dce07bf05d,
64'h9317fdb24face3f8,64'h8fa32e1544e88614,64'h54c740c6eea159d5,64'hffffffff00000000,
64'hc25fa0108f3b0d47,64'h37bc0e9c6b9f4ab0,64'hc6505292cd74e90b,64'h3d212e8cbc8a1ed3,
64'hf40265158762db5d,64'ha5630f77c1b6f3d3,64'hb42cd820857456a5,64'hfffffdff02000201,
64'h537757203e2a1022,64'h054ea8dde9bcdf46,64'hc2aa89fb6115650b,64'hfa4a4eea03df82e5,
64'h98bfed967d671fbc,64'h7d1970ae2744309c,64'ha63a0639750acea6,64'hfffffffefffffff9,
64'h12fd008a79d86a32,64'hbde074e45cfa557f,64'h3282949c6ba74852,64'he9097466e450f697,
64'ha01328b33b16dae1,64'h2b187bc30db79e93,64'ha166c1092ba2b523,64'hffffefff10001001,
64'h9bbab903f150810e,64'h2a7546ef4de6fa30,64'h15544fe108ab2852,64'hd25277571efc1721,
64'hc5ff6cb7eb38fddc,64'he8cb85743a2184dd,64'h31d031d0a856752b,64'hfffffffeffffffc1,
64'h97e80453cec35190,64'hef03a727e7d2abf3,64'h9414a4e45d3a428f,64'h484ba33e2287b4b1,
64'h0099459ed8b6d703,64'h58c3de196dbcf497,64'h0b36084e5d15a913,64'hffff7fff80008001,
64'hddd5c8238a84086c,64'h53aa377b6f37d17f,64'haaa27f0845594290,64'h9293babef7e0b902,
64'h2ffb65c559c7eeda,64'h465c2ba8d10c26e1,64'h8e818e8642b3a957,64'hfffffffefffffe01,
64'hbf4022a2761a8c7c,64'h781d39463e955f91,64'ha0a52726e9d21474,64'h425d19f3143da586,
64'h04ca2cf6c5b6b818,64'hc61ef0cd6de7a4b6,64'h59b04272e8ad4898,64'hfffc000300040001,
64'heeae41225420435a,64'h9d51bbdd79be8bf6,64'h5513f8472aca147b,64'h949dd5fbbf05c80c,
64'h7fdb2e2bce3f76cf,64'h32e15d4888613706,64'h740c7436159d4ab4,64'hfffffffefffff001,
64'hfa011518b0d463db,64'hc0e9ca34f4aafc85,64'h0529393c4e90a39b,64'h12e8cf9aa1ed2c2e,
64'h265167b62db5c0c0,64'h30f786716f3d25aa,64'hcd821399456a44be,64'hffe0001f00200001,
64'h75720919a1021ac9,64'hea8ddeefcdf45fac,64'ha89fc23b5650a3d6,64'ha4eeafe1f82e405c,
64'hfed9716171fbb675,64'h970aea454309b82f,64'ha063a1b3acea559d,64'hfffffffeffff8001,
64'hd008a8cc86a31ed1,64'h074e51ada557e422,64'h2949c9e274851cd8,64'h97467cd50f696170,
64'h328b3db26dae05ff,64'h87bc338c79e92d4f,64'h6c109cd02b5225ea,64'hff0000ff01000001,
64'hab9048d00810d645,64'h546ef7856fa2fd59,64'h44fe11dfb2851eab,64'h27757f14c17202db,
64'hf6cb8b128fddb3a1,64'hb857522e184dc174,64'h031d0da26752ace3,64'hfffffffefffc0001,
64'h8045466a3518f682,64'h3a728d6d2abf2110,64'h4a4e4f14a428e6bf,64'hba33e6ac7b4b0b7c,
64'h9459ed946d702ff7,64'h3de19c67cf496a74,64'h6084e6845a912f4d,64'hf80007ff08000001,
64'h5c8246854086b223,64'ha377bc2d7d17eac6,64'h27f08eff9428f556,64'h3babf8a70b9016d7,
64'hb65c589b7eed9d01,64'hc2ba9175c26e0b9b,64'h18e86d133a956718,64'hfffffffeffe00001,
64'h022a3355a8c7b40c,64'hd3946b6a55f9087f,64'h527278a7214735f6,64'hd19f3568da585bdb,
64'ha2cf6ca76b817fb4,64'hef0ce33f7a4b539f,64'h04273425d4897a65,64'hc0003fff40000001,
64'he412342c04359116,64'h1bbde170e8bf562b,64'h3f8477fda147aaaf,64'hdd5fc5395c80b6b7,
64'hb2e2c4e0f76ce803,64'h15d48bb413705cd2,64'hc7436899d4ab38c0,64'hfffffffeff000001,
64'h11519aad463da060,64'h9ca35b58afc843f2,64'h9393c53b0a39afae,64'h8cf9ab4cd2c2ded2,
64'h167b65405c0bfd9b,64'h78671a02d25a9cf1,64'h2139a12ea44bd328,64'h0002000000000002,
64'h2091a16721ac88a9,64'hddef0b8745fab158,64'hfc23bfee0a3d5577,64'heafe29d0e405b5b2,
64'h9716270cbb674013,64'haea45da09b82e690,64'h3a1b44d4a559c5fa,64'hfffffffef8000001,
64'h8a8cd56a31ed0300,64'he51adac97e421f8c,64'h9c9e29dc51cd7d6c,64'h67cd5a6a9616f68c,
64'hb3db2a02e05fecd8,64'hc338d01992d4e785,64'h09cd0976225e993f,64'h0010000000000010,
64'h048d0b3a0d644547,64'hef785c402fd58aba,64'he11dff7751eaabb1,64'h57f14e8e202dad89,
64'hb8b13869db3a0094,64'h7522ed09dc17347b,64'hd0da26a62ace2fcf,64'hfffffffec0000001,
64'h5466ab558f6817fc,64'h28d6d652f210fc59,64'he4f14ee68e6beb5c,64'h3e6ad357b0b7b45d,
64'h9ed9501c02ff66bb,64'h19c680d296a73c22,64'h4e684bb112f4c9f8,64'h0080000000000080,
64'h246859d06b222a38,64'h7bc2e2087eac55c9,64'h08effbc18f555d81,64'hbf8a7473016d6c46,
64'hc589c353d9d0049b,64'ha9176851e0b9a3d5,64'h86d1353756717e72,64'hfffffffd00000001,
64'ha3355aae7b40bfde,64'h46b6b2989087e2c7,64'h278a773b735f5ad9,64'hf3569abe85bda2e7,
64'hf6ca80e417fb35d4,64'hce340694b539e110,64'h73425d8a97a64fbe,64'h0400000000000400,
64'h2342ce84591151bf,64'hde171046f562ae45,64'h477fde0c7aaaec08,64'hfc53a39d0b6b622b,
64'h2c4e1aa4ce8024d2,64'h48bb429405cd1ea3,64'h3689a9beb38bf38c,64'hffffffef00000001,
64'h19aad578da05feeb,64'h35b594c6843f1636,64'h3c53b9dc9afad6c7,64'h9ab4d5fb2ded1731,
64'hb6540727bfd9ae99,64'h71a034aba9cf087a,64'h9a12ec57bd327ded,64'h2000000000002000,
64'h1a167423c88a8df7,64'hf0b8823dab157222,64'h3bfef065d557603e,64'he29d1cef5b5b1151,
64'h6270d5277401268f,64'h45da14a22e68f516,64'hb44d4df69c5f9c5f,64'hffffff7f00000001,
64'hcd56abc6d02ff758,64'hadaca63521f8b1af,64'he29dcee5d7d6b637,64'hd5a6afdd6f68b984,
64'hb2a03942fecd74c3,64'h8d01a5604e7843cd,64'hd09762c1e993ef64,64'h000000010000ffff,
64'hd0b3a11e44546fb8,64'h85c411f458ab9109,64'hdff7832faabb01ef,64'h14e8e781dad88a81,
64'h1386a93ea0093475,64'h2ed0a5137347a8ae,64'ha26a6fb9e2fce2f3,64'hfffffbff00000001,
64'h6ab55e3c817fbaba,64'h6d6531ae0fc58d73,64'h14ee7735beb5b1b1,64'had357ef17b45cc1a,
64'h9501ca1cf66ba613,64'h680d2b0673c21e64,64'h84bb16154c9f7b1a,64'h000000080007fff8,
64'h859d08f822a37dba,64'h2e208fa6c55c8844,64'hffbc198355d80f72,64'ha7473c0ed6c45408,
64'h9c3549f50049a3a8,64'h7685289c9a3d456f,64'h13537dd417e71793,64'hffffdfff00000001,
64'h55aaf1e70bfdd5cd,64'h6b298d737e2c6b95,64'ha773b9adf5ad8d88,64'h69abf790da2e60cb,
64'ha80e50ebb35d3094,64'h406958369e10f31d,64'h25d8b0ae64fbd8cc,64'h00000040003fffc0,
64'h2ce847c5151bedcc,64'h71047d372ae4421f,64'hfde0cc21aec07b89,64'h3a39e07bb622a03b,
64'he1aa4fac024d1d3c,64'hb42944e7d1ea2b75,64'h9a9beea0bf38bc98,64'hfffeffff00000001,
64'had578f3a5feeae66,64'h594c6b9ef1635ca5,64'h3b9dcd74ad6c6c3b,64'h4d5fbc89d1730655,
64'h407287629ae9849b,64'h034ac1b6f08798e6,64'h2ec5857427dec65f,64'h0000020001fffe00,
64'h67423e29a8df6e5f,64'h8823e9bc572210f5,64'hef0661147603dc41,64'hd1cf03deb11501d7,
64'h0d527d671268e9d9,64'ha14a27438f515ba3,64'hd4df7509f9c5e4bc,64'hfff7ffff00000001,
64'h6abc79d7ff75732b,64'hca635cf98b1ae526,64'hdcee6ba66b6361d7,64'h6afde4508b9832a6,
64'h03943b16d74c24d6,64'h1a560db7843cc730,64'h762c2ba23ef632f7,64'h000010000ffff000,
64'h3a11f15046fb72f5,64'h411f4de6b91087a4,64'h783308aab01ee201,64'h8e781efb88a80eb2,
64'h6a93eb3893474ec8,64'h0a513a217a8add13,64'ha6fba855ce2f25da,64'hffbfffff00000001,
64'h55e3cec2fbab9955,64'h531ae7d258d7292a,64'he7735d395b1b0eb2,64'h57ef22875cc1952d,
64'h1ca1d8b6ba6126b0,64'hd2b06dbc21e63980,64'hb1615d14f7b197b5,64'h000080007fff8000,
64'hd08f8a8337db97a7,64'h08fa6f37c8843d1e,64'hc198455880f71005,64'h73c0f7e04540758c,
64'h549f59c79a3a763d,64'h5289d10bd456e898,64'h37dd42b371792ecb,64'hfdffffff00000001,
64'haf1e7619dd5ccaa6,64'h98d73e94c6b9494e,64'h3b9ae9d1d8d87589,64'hbf79143ce60ca966,
64'he50ec5b5d3093580,64'h95836de70f31cbfa,64'h8b0ae8acbd8cbda3,64'h00040003fffc0000,
64'h847c541fbedcbd32,64'h47d379be4421e8f0,64'h0cc22aca07b88022,64'h9e07bf052a03ac5d,
64'ha4face3ed1d3b1e6,64'h944e8860a2b744be,64'hbeea159c8bc97657,64'hefffffff00000001,
64'h78f3b0d3eae6552b,64'hc6b9f4aa35ca4a6c,64'hdcd74e8fc6c3ac47,64'hfbc8a1ec30654b2b,
64'h28762db59849abf9,64'hac1b6f3c798e5fcc,64'h58574569ec65ed14,64'h0020001fffe00000,
64'h23e2a101f6e5e98c,64'h3e9bcdf4210f477e,64'h661156503dc40110,64'hf03df82d501d62e4,
64'h27d671fb8e9d8f2b,64'ha274430915ba25ec,64'hf750ace95e4bb2b3,64'h7fffffff00000001,
64'hc79d86a25732a955,64'h35cfa557ae52535a,64'he6ba7484361d6232,64'hde450f68832a5951,
64'h43b16dadc24d5fc7,64'h60db79e8cc72fe5b,64'hc2ba2b51632f689e,64'h010000ffff000000,
64'h1f150810b72f4c5f,64'hf4de6fa2087a3bef,64'h308ab284ee20087d,64'h81efc17180eb1719,
64'h3eb38fdd74ec7957,64'h13a2184dadd12f5b,64'hba856751f25d9591,64'hfffffffb00000005,
64'h3cec3518b9954aa2,64'hae7d2abe72929acf,64'h35d3a428b0eb1189,64'hf2287b4a1952ca82,
64'h1d8b6d70126afe36,64'h06dbcf496397f2d5,64'h15d15a91197b44ea,64'h080007fff8000000,
64'hf8a84085b97a62f8,64'ha6f37d1743d1df71,64'h84559428710043e7,64'h0f7e0b900758b8c4,
64'hf59c7eeca763cab7,64'h9d10c26d6e897ad8,64'hd42b3a9492ecac83,64'hffffffdf00000021,
64'he761a8c6ccaa550f,64'h73e955f89494d673,64'hae9d214687588c47,64'h9143da57ca965409,
64'hec5b6b809357f1b0,64'h36de7a4b1cbf96a8,64'hae8ad488cbda2750,64'h40003fffc0000000,
64'hc5420434cbd317b9,64'h379be8bf1e8efb83,64'h22aca14788021f34,64'h7bf05c803ac5c620,
64'hace3f76c3b1e55b1,64'he886136f744bd6bc,64'ha159d4aa97656412,64'hfffffeff00000101,
64'h3b0d463d6552a871,64'h9f4aafc7a4a6b395,64'h74e90a393ac46233,64'h8a1ed2c254b2a044,
64'h62db5c0b9abf8d79,64'hb6f3d259e5fcb53f,64'h7456a44b5ed13a7b,64'h0001fffffffffffe,
64'h2a1021ac5e98bdc2,64'hbcdf45f9f477dc17,64'h15650a3d4010f99f,64'hdf82e404d62e30fd,
64'h671fbb66d8f2ad83,64'h44309b82a25eb5d9,64'h0acea559bb2b208b,64'hfffff7ff00000801,
64'hd86a31ec2a954387,64'hfa557e4125359ca4,64'ha74851ccd6231195,64'h50f69616a595021c,
64'h16dae05fd5fc6bc5,64'hb79e92d42fe5a9f3,64'ha2b5225df689d3d5,64'h000ffffffffffff0,
64'h50810d63f4c5ee0f,64'he6fa2fd4a3bee0b3,64'hab2851ea0087ccf8,64'hfc17202cb17187e2,
64'h38fddb39c7956c15,64'h2184dc1712f5aec6,64'h56752acdd9590458,64'hffffbfff00004001,
64'hc3518f6754aa1c32,64'hd2abf21029ace519,64'h3a428e6bb1188ca3,64'h87b4b0b72ca810de,
64'hb6d702feafe35e28,64'hbcf496a67f2d4f93,64'h15a912f4b44e9ea3,64'h007fffffffffff80,
64'h84086b21a62f7076,64'h37d17eac1df70591,64'h59428f55043e67bb,64'he0b9016c8b8c3f09,
64'hc7eed9cf3cab60a7,64'h0c26e0b997ad762f,64'hb3a95670cac822be,64'hfffdffff00020001,
64'h1a8c7b40a550e18a,64'h955f90874d6728c2,64'hd214735e88c46517,64'h3da585bd654086ec,
64'hb6b817fa7f1af13b,64'he7a4b538f96a7c93,64'had4897a5a274f518,64'h03fffffffffffc00,
64'h20435911317b83ac,64'hbe8bf561efb82c87,64'hca147aaa21f33dd6,64'h05c80b6b5c61f841,
64'h3f76ce7fe55b0532,64'h613705ccbd6bb178,64'h9d4ab38b564115eb,64'hffefffff00100001,
64'hd463da052a870c50,64'haafc843e6b39460c,64'h90a39afa462328b2,64'hed2c2dec2a04375f,
64'hb5c0bfd8f8d789d3,64'h3d25a9cecb53e491,64'h6a44bd3213a7a8bb,64'h1fffffffffffe000,
64'h021ac88a8bdc1d5f,64'hf45fab147dc16433,64'h50a3d5570f99eeaa,64'h2e405b5ae30fc208,
64'hfbb674002ad8298f,64'h09b82e68eb5d8bbd,64'hea559c5eb208af54,64'hff7fffff00800001
};
  //------------------------
  // 256
  //------------------------
  localparam [2*256-1:0][63:0] NTT_GF64_BWD_WDIV_N256_PHI_L = {
64'hafc843f0b39460b6,64'hd2c2ded0a04375e2,64'hd25a9cefb53e490d,64'h00000001fffdfffe,
64'h45fab156dc164321,64'he405b5b030fc207e,64'h9b82e68eb5d8bbd0,64'hf7ffffff08000001,
64'h7e421f8a9ca305ab,64'h9616f68b021baf0a,64'h92d4e783a9f24862,64'h0000000fffeffff0,
64'h2fd58ab8e0b21906,64'h202dad8887e103e9,64'hdc173479aec5de7c,64'hbfffffff40000001,
64'hf210fc57e5182d55,64'hb0b7b45c10dd784c,64'h96a73c214f92430c,64'h0000007fff7fff80,
64'h7eac55c80590c82f,64'h016d6c453f081f47,64'he0b9a3d3762ef3da,64'h0000000000000002,
64'h9087e2c628c16aa1,64'h85bda2e586ebc25b,64'hb539e10e7c92185c,64'h000003fffbfffc00,
64'hf562ae432c864175,64'h0b6b6229f840fa38,64'h05cd1ea2b1779ec9,64'h0000000000000010,
64'h843f1635460b5504,64'h2ded1730375e12d4,64'ha9cf0878e490c2db,64'h00001fffdfffe000,
64'hab15722064320ba1,64'h5b5b114fc207d1c0,64'h2e68f5158bbcf648,64'h0000000000000080,
64'h21f8b1ae305aa81c,64'h6f68b982baf0969f,64'h4e7843cc248616d3,64'h0000fffeffff0000,
64'h58ab910821905d03,64'hdad88a80103e8dfe,64'h7347a8ad5de7b23f,64'h0000000000000400,
64'h0fc58d7282d540df,64'h7b45cc18d784b4f5,64'h73c21e632430b696,64'h0007fff7fff80000,
64'hc55c88430c82e816,64'hd6c4540681f46fea,64'h9a3d456def3d91f5,64'h0000000000002000,
64'h7e2c6b9416aa06f8,64'hda2e60c9bc25a7a5,64'h9e10f31c2185b4ad,64'h003fffbfffc00000,
64'h2ae4421e641740aa,64'hb622a03a0fa37f4a,64'hd1ea2b7379ec8fa4,64'h0000000000010000,
64'hf1635ca3b55037bd,64'hd1730653e12d3d22,64'hf08798e50c2da564,64'h01fffdfffe000000,
64'h572210f420ba054f,64'hb11501d57d1bfa4b,64'h8f515ba1cf647d1a,64'h0000000000080000,
64'h8b1ae524aa81bde1,64'h8b9832a50969e90a,64'h843cc72f616d2b19,64'h0fffeffff0000000,
64'hb91087a305d02a76,64'h88a80eb0e8dfd253,64'h7a8add127b23e8cc,64'h0000000000400000,
64'h58d72929540def04,64'h5cc1952c4b4f484c,64'h21e6397f0b6958c4,64'h7fff7fff80000000,
64'hc8843d1d2e8153ab,64'h4540758b46fe9294,64'hd456e896d91f465d,64'h0000000002000000,
64'hc6b9494ca06f781e,64'he60ca9645a7a425e,64'h0f31cbf95b4ac61f,64'hfffbfffefffffffd,
64'h4421e8ef740a9d52,64'h2a03ac5c37f4949e,64'ha2b744bcc8fa32e2,64'h0000000010000000,
64'h35ca4a6b037bc0ea,64'h30654b29d3d212e9,64'h798e5fcada5630f8,64'hffdffffeffffffe1,
64'h210f477da054ea8e,64'h501d62e2bfa4a4ef,64'h15ba25eb47d1970b,64'h0000000080000000,
64'hae5253591bde074f,64'h832a594f9e909747,64'hcc72fe59d2b187bd,64'hfefffffeffffff01,
64'h087a3bee02a7546f,64'h80eb1717fd252776,64'hadd12f5a3e8cb858,64'h0000000400000000,
64'h72929acddef03a73,64'h1952ca80f484ba34,64'h6397f2d4958c3de2,64'hf7fffffefffff801,
64'h43d1df70153aa378,64'h0758b8c3e9293bac,64'h6e897ad6f465c2bb,64'h0000002000000000,
64'h9494d671f781d395,64'hca965407a425d1a0,64'h1cbf96a7ac61ef0d,64'hbffffffeffffc001,
64'h1e8efb82a9d51bbe,64'h3ac5c61f4949dd60,64'h744bd6baa32e15d5,64'h0000010000000000,
64'ha4a6b393bc0e9ca4,64'h54b2a043212e8cfa,64'he5fcb53d630f7868,64'hfffffffcfffe0003,
64'hf477dc154ea8ddf0,64'hd62e30fb4a4eeaff,64'ha25eb5d81970aea5,64'h0000080000000000,
64'h25359ca2e074e51b,64'ha595021b097467ce,64'h2fe5a9f2187bc339,64'hffffffeefff00011,
64'ha3bee0b17546ef79,64'hb17187e0527757f2,64'h12f5aec5cb857523,64'h0000400000000000,
64'h29ace51803a728d7,64'h2ca810dd4ba33e6b,64'h7f2d4f91c3de19c7,64'hffffff7eff800081,
64'h1df70590aa377bc3,64'h8b8c3f0793babf8b,64'h97ad762e5c2ba918,64'h0002000000000000,
64'h4d6728c11d3946b7,64'h654086eb5d19f357,64'hf96a7c911ef0ce35,64'hfffffbfefc000401,
64'hefb82c8551bbde18,64'h5c61f8409dd5fc54,64'hbd6bb176e15d48bc,64'h0010000000000000,
64'h6b39460ae9ca35b6,64'h2a04375de8cf9ab5,64'hcb53e48ff78671a1,64'hffffdffee0002001,
64'h7dc164318ddef0b9,64'he30fc206eeafe29e,64'heb5d8bbc0aea45db,64'h0080000000000000,
64'h59ca305a4e51adad,64'h5021baf0467cd5a7,64'h5a9f2485bc338d02,64'hfffefffe00010001,
64'hee0b218f6ef785c5,64'h187e103e757f14e9,64'h5aec5de757522ed1,64'h0400000000000000,
64'hce5182d4728d6d66,64'h810dd78433e6ad36,64'hd4f9242fe19c680e,64'hfff7fff700080001,
64'h70590c8277bc2e21,64'hc3f081f3abf8a748,64'hd762ef3cba917686,64'h2000000000000000,
64'h728c16a9946b6b2a,64'h086ebc259f3569ac,64'ha7c921850ce3406a,64'hffbfffbf00400001,
64'h82c86416bde17105,64'h1f840fa35fc53a3a,64'hbb1779ebd48bb42a,64'h00000000ffffffff,
64'h9460b54fa35b594d,64'h4375e12cf9ab4d60,64'h3e490c2d671a034b,64'hfdfffdff02000001,
64'h164320b9ef0b8824,64'hfc207d1afe29d1d0,64'hd8bbcf63a45da14b,64'h00000007fffffff8,
64'ha305aa811adaca64,64'h1baf0969cd5a6afe,64'hf248616c38d01a57,64'hefffefff10000001,
64'hb21905cf785c4120,64'he103e8def14e8e79,64'hc5de7b2322ed0a52,64'h0000003fffffffc0,
64'h182d540dd6d6531b,64'hdd784b4e6ad357f0,64'h92430b68c680d2b1,64'h7fff7fff80000001,
64'h90c82e80c2e208fb,64'h081f46fe8a7473c1,64'h2ef3d91f1768528a,64'h000001fffffffe00,
64'hc16aa06eb6b298d8,64'hebc25a79569abf7a,64'h92185b4a34069584,64'hfffbffff00000005,
64'h8641740a171047d4,64'h40fa37f453a39e08,64'h779ec8f9bb42944f,64'h00000ffffffff000,
64'h0b55037bb594c6ba,64'h5e12d3d1b4d5fbc9,64'h90c2da55a034ac1c,64'hffdfffff00000021,
64'h320ba054b8823e9c,64'h07d1bfa49d1cf03e,64'hbcf647d0da14a275,64'h00007fffffff8000,
64'h5aa81bddaca635d0,64'hf0969e8fa6afde46,64'h8616d2b101a560dc,64'hfeffffff00000101,
64'h905d02a6c411f4df,64'h3e8dfd24e8e781f0,64'he7b23e8bd0a513a3,64'h0003fffffffc0000,
64'hd540deef6531ae7e,64'h84b4f484357ef229,64'h30b6958c0d2b06dc,64'hf7ffffff00000801,
64'h82e8153a208fa6f4,64'hf46fe928473c0f7f,64'h3d91f46585289d11,64'h001fffffffe00000,
64'haa06f781298d73ea,64'h25a7a425abf79144,64'h85b4ac61695836df,64'hbfffffff00004001,
64'h1740a9d5047d379c,64'ha37f494939e07bf1,64'hec8fa32d2944e887,64'h00ffffffff000000,
64'h5037bc0e4c6b9f4b,64'h2d3d212e5fbc8a1f,64'h2da5630f4ac1b6f4,64'hfffffffd00020003,
64'hba054ea823e9bce0,64'h1bfa4a4ecf03df83,64'h647d19704a274431,64'h07fffffff8000000,
64'h81bde074635cfa56,64'h69e90973fde450f7,64'h6d2b187b560db79f,64'hffffffef00100011,
64'hd02a75461f4de6fb,64'hdfd25276781efc18,64'h23e8cb85513a2185,64'h3fffffffc0000000,
64'h0def03a71ae7d2ac,64'h4f484ba2ef2287b5,64'h6958c3ddb06dbcf5,64'hffffff7f00800081,
64'h8153aa36fa6f37d2,64'hfe9293b9c0f7e0ba,64'h1f465c2b89d10c27,64'hfffffffeffffffff,
64'h6f781d38d73e9560,64'h7a425d1979143da6,64'h4ac61ef0836de7a5,64'hfffffbff04000401,
64'h0a9d51bbd379be8c,64'hf4949dd507bf05c9,64'hfa32e15c4e886138,64'hfffffffefffffff1,
64'h7bc0e9c9b9f4aafd,64'hd212e8cec8a1ed2d,64'h5630f7861b6f3d26,64'hffffdfff20002001,
64'h54ea8dde9bcdf460,64'ha4a4eeaf3df82e41,64'hd1970ae9744309b9,64'hfffffffeffffff81,
64'hde074e50cfa557e5,64'h9097467c450f6962,64'hb187bc32db79e92e,64'hffff000000010001,
64'ha7546ef6de6fa2fe,64'h2527757eefc17203,64'h8cb85751a2184dc2,64'hfffffffefffffc01,
64'hf03a728c7d2abf22,64'h84ba33e6287b4b0c,64'h8c3de19bdbcf496b,64'hfff8000700080001,
64'h3aa377bbf37d17eb,64'h293babf87e0b9017,64'h65c2ba9110c26e0c,64'hfffffffeffffe001,
64'h81d3946ae955f909,64'h25d19f3543da585c,64'h61ef0ce2de7a4b54,64'hffc0003f00400001,
64'hd51bbde09be8bf57,64'h49dd5fc4f05c80b7,64'h2e15d48b8613705d,64'hfffffffeffff0001,
64'h0e9ca35b4aafc844,64'h2e8cf9ab1ed2c2df,64'h0f786719f3d25a9d,64'hfe0001ff02000001,
64'ha8ddef0adf45fab2,64'h4eeafe2982e405b6,64'h70aea45d309b82e7,64'hfffffffefff80001,
64'h74e51ada557e4220,64'h7467cd59f69616f7,64'h7bc338cf9e92d4e8,64'hf0000fff10000001,
64'h46ef785bfa2fd58b,64'h7757f14e17202dae,64'h857522ec84dc1735,64'hfffffffeffc00001,
64'ha728d6d5abf210fd,64'ha33e6ad2b4b0b7b5,64'hde19c67ff496a73d,64'h80007fff80000001,
64'h377bc2e1d17eac56,64'hbabf8a73b9016d6d,64'h2ba9176826e0b9a4,64'hfffffffefe000001,
64'h3946b6b25f9087e3,64'h19f3569aa585bda3,64'hf0ce3405a4b539e2,64'h0004000000000004,
64'hbbde170f8bf562af,64'hd5fc53a2c80b6b63,64'h5d48bb423705cd1f,64'hfffffffef0000001,
64'hca35b593fc843f17,64'hcf9ab4d52c2ded18,64'h8671a03425a9cf09,64'h0020000000000020,
64'hdef0b8815fab1573,64'hafe29d1c405b5b12,64'hea45da13b82e68f6,64'hfffffffe80000001,
64'h51adaca5e421f8b2,64'h7cd5a6af616f68ba,64'h338d01a52d4e7844,64'h0100000000000100,
64'hf785c410fd58ab92,64'h7f14e8e702dad88b,64'h522ed0a4c17347a9,64'hfffffffb00000001,
64'h8d6d6531210fc58e,64'he6ad357e0b7b45cd,64'h9c680d2a6a73c21f,64'h0800000000000800,
64'hbc2e208eeac55c89,64'hf8a7473b16d6c455,64'h917685280b9a3d46,64'hffffffdf00000001,
64'h6b6b298d087e2c6c,64'h3569abf75bda2e61,64'he3406957539e10f4,64'h4000000000004000,
64'he171047c562ae443,64'hc53a39dfb6b622a1,64'h8bb429445cd1ea2c,64'hfffffeff00000001,
64'h5b594c6b43f1635d,64'hab4d5fbbded17307,64'h1a034ac19cf08799,64'h000000020001fffe,
64'h0b8823e9b1572211,64'h29d1cf03b5b11502,64'h5da14a26e68f515c,64'hfffff7ff00000001,
64'hdaca635c1f8b1ae6,64'h5a6afde3f68b9833,64'hd01a560ce7843cc8,64'h00000010000ffff0,
64'h5c411f4d8ab91088,64'h4e8e781ead88a80f,64'hed0a5139347a8ade,64'hffffbfff00000001,
64'hd6531ae6fc58d72a,64'hd357ef21b45cc196,64'h80d2b06d3c21e63a,64'h00000080007fff80,
64'he208fa6e55c8843e,64'h7473c0f76c454076,64'h685289d0a3d456e9,64'hfffdffff00000001,
64'hb298d73de2c6b94a,64'h9abf7913a2e60caa,64'h0695836de10f31cc,64'h0000040003fffc00,
64'h1047d379ae4421e9,64'ha39e07be622a03ad,64'h42944e881ea2b745,64'hffefffff00000001,
64'h94c6b9f41635ca4b,64'hd5fbc8a11730654c,64'h34ac1b6f08798e60,64'h000020001fffe000,
64'h823e9bcd72210f48,64'h1cf03df811501d63,64'h14a27442f515ba26,64'hff7fffff00000001,
64'ha635cfa4b1ae5254,64'hafde450eb9832a5a,64'ha560db7943cc72ff,64'h00010000ffff0000,
64'h11f4de6f91087a3c,64'he781efc08a80eb18,64'ha513a217a8add130,64'hfbffffff00000001,
64'h31ae7d2a8d72929b,64'h7ef2287acc1952cb,64'h2b06dbcf1e6397f3,64'h00080007fff80000,
64'h8fa6f37c8843d1e0,64'h3c0f7e0b540758b9,64'h289d10c2456e897b,64'hdfffffff00000001,
64'h8d73e9556b9494d7,64'hf79143d960ca9655,64'h5836de79f31cbf97,64'h0040003fffc00000,
64'h7d379be8421e8efc,64'he07bf05ba03ac5c7,64'h44e886132b744bd7,64'hfffffffe00000002,
64'h6b9f4aaf5ca4a6b4,64'hbc8a1ed20654b2a1,64'hc1b6f3d198e5fcb6,64'h020001fffe000000,
64'he9bcdf4510f477dd,64'h03df82e401d62e31,64'h2744309b5ba25eb6,64'hfffffff700000009,
64'h5cfa557de525359d,64'he450f69532a59503,64'h0db79e92c72fe5aa,64'h10000ffff0000000,
64'h4de6fa2f87a3bee1,64'h1efc17200eb17188,64'h3a2184dbdd12f5af,64'hffffffbf00000041,
64'he7d2abf12929ace6,64'h2287b4b0952ca811,64'h6dbcf496397f2d50,64'h80007fff80000000,
64'h6f37d17e3d1df706,64'hf7e0b900758b8c40,64'hd10c26dfe897ad77,64'hfffffdff00000201,
64'h3e955f90494d6729,64'h143da585a9654087,64'h6de7a4b4cbf96a7d,64'h0003fffffffffffc,
64'h79be8bf4e8efb82d,64'hbf05c80aac5c61f9,64'h8861370544bd6bb2,64'hffffefff00001001,
64'hf4aafc834a6b3947,64'ha1ed2c2d4b2a0438,64'h6f3d25a95fcb53e5,64'h001fffffffffffe0,
64'hcdf45faa477dc165,64'hf82e405a62e30fc3,64'h4309b82e25eb5d8c,64'hffff7fff00008001,
64'ha557e4215359ca31,64'h0f69616f595021bb,64'h79e92d4dfe5a9f25,64'h00ffffffffffff00,
64'h6fa2fd583bee0b22,64'hc17202da17187e11,64'h184dc1732f5aec5e,64'hfffbffff00040001,
64'h2abf210f9ace5183,64'h7b4b0b7aca810dd8,64'hcf496a72f2d4f925,64'h07fffffffffff800,
64'h7d17eac4df70590d,64'h0b9016d6b8c3f082,64'hc26e0b997ad762f0,64'hffdfffff00200001,
64'h55f9087dd6728c17,64'hda585bd954086ebd,64'h7a4b539d96a7c922,64'h3fffffffffffc000,
64'he8bf5629fb82c865,64'h5c80b6b5c61f8410,64'h13705cd1d6bb177a,64'hfeffffff01000001
};
  //------------------------
  // 128
  //------------------------
  localparam [2*128-1:0][63:0] NTT_GF64_BWD_WDIV_N128_PHI_L = {
64'ha585bda24086ebc3,64'h00000003fffbfffc,64'hc80b6b6161f840fb,64'hefffffff10000001,
64'h2c2ded1704375e13,64'h0000001fffdfffe0,64'h405b5b110fc207d2,64'h7fffffff80000001,
64'h616f68b921baf097,64'h000000fffeffff00,64'h02dad88a7e103e8e,64'h0000000000000004,
64'h0b7b45cc0dd784b5,64'h000007fff7fff800,64'h16d6c453f081f470,64'h0000000000000020,
64'h5bda2e606ebc25a8,64'h00003fffbfffc000,64'hb6b6229f840fa380,64'h0000000000000100,
64'hded1730575e12d3e,64'h0001fffdfffe0000,64'hb5b11501207d1bfb,64'h0000000000000800,
64'hf68b9831af0969ea,64'h000fffeffff00000,64'had88a80e03e8dfd3,64'h0000000000004000,
64'hb45cc194784b4f49,64'h007fff7fff800000,64'h6c4540751f46fe93,64'h0000000000020000,
64'ha2e60ca8c25a7a43,64'h03fffbfffc000000,64'h622a03abfa37f495,64'h0000000000100000,
64'h1730654b12d3d213,64'h1fffdfffe0000000,64'h11501d62d1bfa4a5,64'h0000000000800000,
64'hb9832a58969e9098,64'hfffeffff00000000,64'h8a80eb168dfd2528,64'h0000000004000000,
64'hcc1952c9b4f484bb,64'hfff7fffefffffff9,64'h540758b86fe9293c,64'h0000000020000000,
64'h60ca9653a7a425d2,64'hffbffffeffffffc1,64'ha03ac5c57f4949de,64'h0000000100000000,
64'h0654b2a03d212e8d,64'hfdfffffefffffe01,64'h01d62e30fa4a4eeb,64'h0000000800000000,
64'h32a59501e9097468,64'heffffffefffff001,64'h0eb17187d2527758,64'h0000004000000000,
64'h952ca810484ba33f,64'h7ffffffeffff8001,64'h758b8c3e9293bac0,64'h0000020000000000,
64'ha9654086425d19f4,64'hfffffffafffc0005,64'hac5c61f7949dd5fd,64'h0000100000000000,
64'h4b2a043712e8cf9b,64'hffffffdeffe00021,64'h62e30fc1a4eeafe3,64'h0000800000000000,
64'h595021ba97467cd6,64'hfffffefeff000101,64'h17187e1027757f15,64'h0004000000000000,
64'hca810dd6ba33e6ae,64'hfffff7fef8000801,64'hb8c3f0813babf8a8,64'h0020000000000000,
64'h54086ebbd19f356a,64'hffffbffec0004001,64'hc61f840edd5fc53b,64'h0100000000000000,
64'ha04375e08cf9ab4e,64'hfffdfffd00020001,64'h30fc207ceafe29d2,64'h0800000000000000,
64'h021baf0967cd5a6b,64'hffefffef00100001,64'h87e103e857f14e8f,64'h4000000000000000,
64'h10dd784b3e6ad358,64'hff7fff7f00800001,64'h3f081f46bf8a7474,64'h00000001fffffffe,
64'h86ebc259f3569ac0,64'hfbfffbff04000001,64'hf840fa36fc53a39f,64'h0000000ffffffff0,
64'h375e12d39ab4d5fc,64'hdfffdfff20000001,64'hc207d1bee29d1cf1,64'h0000007fffffff80,
64'hbaf0969dd5a6afdf,64'hfffeffff00000002,64'h103e8dfd14e8e782,64'h000003fffffffc00,
64'hd784b4f3ad357ef3,64'hfff7ffff00000009,64'h81f46fe8a7473c10,64'h00001fffffffe000,
64'hbc25a7a369abf792,64'hffbfffff00000041,64'h0fa37f493a39e07c,64'h0000ffffffff0000,
64'he12d3d204d5fbc8b,64'hfdffffff00000201,64'h7d1bfa49d1cf03e0,64'h0007fffffff80000,
64'h0969e9096afde451,64'hefffffff00001001,64'he8dfd2518e781efd,64'h003fffffffc00000,
64'h4b4f484b57ef2288,64'h7fffffff00008001,64'h46fe929373c0f7e1,64'h01fffffffe000000,
64'h5a7a425cbf79143e,64'hfffffffb00040005,64'h37f4949d9e07bf06,64'h0ffffffff0000000,
64'hd3d212e7fbc8a1ee,64'hffffffdf00200021,64'hbfa4a4edf03df82f,64'h7fffffff80000000,
64'h9e909745de450f6a,64'hfffffeff01000101,64'hfd25277481efc173,64'hfffffffefffffffd,
64'hf484ba32f2287b4c,64'hfffff7ff08000801,64'he9293bab0f7e0b91,64'hfffffffeffffffe1,
64'ha425d19e9143da59,64'hffffbfff40004001,64'h4949dd5f7bf05c81,64'hfffffffeffffff01,
64'h212e8cf98a1ed2c3,64'hfffe000100020001,64'h4a4eeafddf82e406,64'hfffffffefffff801,
64'h097467cd50f69617,64'hfff0000f00100001,64'h527757f0fc17202e,64'hfffffffeffffc001,
64'h4ba33e6a87b4b0b8,64'hff80007f00800001,64'h93babf89e0b9016e,64'hfffffffefffe0001,
64'h5d19f3563da585be,64'hfc0003ff04000001,64'h9dd5fc5305c80b6c,64'hfffffffefff00001,
64'he8cf9ab3ed2c2dee,64'he0001fff20000001,64'heeafe29c2e405b5c,64'hfffffffeff800001,
64'h467cd5a669616f69,64'h0001000000000001,64'h757f14e87202dad9,64'hfffffffefc000001,
64'h33e6ad354b0b7b46,64'h0008000000000008,64'habf8a7469016d6c5,64'hfffffffee0000001,
64'h9f3569ab585bda2f,64'h0040000000000040,64'h5fc53a3980b6b623,64'hfffffffe00000001,
64'hf9ab4d5ec2ded174,64'h0200000000000200,64'hfe29d1ce05b5b116,64'hfffffff700000001,
64'hcd5a6afd16f68b99,64'h1000000000001000,64'hf14e8e772dad88a9,64'hffffffbf00000001,
64'h6ad357eeb7b45cc2,64'h8000000000008000,64'h8a7473c06d6c4541,64'hfffffdff00000001,
64'h569abf78bda2e60d,64'h000000040003fffc,64'h53a39e076b622a04,64'hffffefff00000001,
64'hb4d5fbc7ed173066,64'h00000020001fffe0,64'h9d1cf03d5b11501e,64'hffff7fff00000001,
64'ha6afde4468b9832b,64'h0000010000ffff00,64'he8e781eed88a80ec,64'hfffbffff00000001,
64'h357ef22845cc1953,64'h0000080007fff800,64'h473c0f7dc4540759,64'hffdfffff00000001,
64'habf791432e60ca97,64'h000040003fffc000,64'h39e07bf022a03ac6,64'hfeffffff00000001,
64'h5fbc8a1e730654b3,64'h00020001fffe0000,64'hcf03df821501d62f,64'hf7ffffff00000001,
64'hfde450f59832a596,64'h0010000ffff00000,64'h781efc16a80eb172,64'hbfffffff00000001,
64'hef2287b3c1952ca9,64'h0080007fff800000,64'hc0f7e0b840758b8d,64'hfffffffd00000003,
64'h79143da50ca96541,64'h040003fffc000000,64'h07bf05c803ac5c62,64'hffffffef00000011,
64'hc8a1ed2b654b2a05,64'h20001fffe0000000,64'h3df82e401d62e310,64'hffffff7f00000081,
64'h450f69612a595022,64'h0000ffffffffffff,64'hefc17201eb17187f,64'hfffffbff00000401,
64'h287b4b0b52ca810e,64'h0007fffffffffff8,64'h7e0b901658b8c3f1,64'hffffdfff00002001,
64'h43da585b9654086f,64'h003fffffffffffc0,64'hf05c80b5c5c61f85,64'hfffeffff00010001,
64'h1ed2c2deb2a04376,64'h01fffffffffffe00,64'h82e405b52e30fc21,64'hfff7ffff00080001,
64'hf69616f595021bb0,64'h0ffffffffffff000,64'h17202dad7187e104,64'hffbfffff00400001,
64'hb4b0b7b3a810dd79,64'h7fffffffffff8000,64'hb9016d6b8c3f0820,64'hfdffffff02000001
};
  //------------------------
  // 64
  //------------------------
  localparam [2*64-1:0][63:0] NTT_GF64_BWD_WDIV_N64_PHI_L = {
64'h00000007fff7fff8,64'hdfffffff20000001,64'h0000003fffbfffc0,64'h0000000000000001,
64'h000001fffdfffe00,64'h0000000000000008,64'h00000fffeffff000,64'h0000000000000040,
64'h00007fff7fff8000,64'h0000000000000200,64'h0003fffbfffc0000,64'h0000000000001000,
64'h001fffdfffe00000,64'h0000000000008000,64'h00fffeffff000000,64'h0000000000040000,
64'h07fff7fff8000000,64'h0000000000200000,64'h3fffbfffc0000000,64'h0000000001000000,
64'hfffdfffeffffffff,64'h0000000008000000,64'hffeffffefffffff1,64'h0000000040000000,
64'hff7ffffeffffff81,64'h0000000200000000,64'hfbfffffefffffc01,64'h0000001000000000,
64'hdffffffeffffe001,64'h0000008000000000,64'hfffffffdffff0002,64'h0000040000000000,
64'hfffffff6fff80009,64'h0000200000000000,64'hffffffbeffc00041,64'h0001000000000000,
64'hfffffdfefe000201,64'h0008000000000000,64'hffffeffef0001001,64'h0040000000000000,
64'hffff7ffe80008001,64'h0200000000000000,64'hfffbfffb00040001,64'h1000000000000000,
64'hffdfffdf00200001,64'h8000000000000000,64'hfefffeff01000001,64'h00000003fffffffc,
64'hf7fff7ff08000001,64'h0000001fffffffe0,64'hbfffbfff40000001,64'h000000ffffffff00,
64'hfffdffff00000003,64'h000007fffffff800,64'hffefffff00000011,64'h00003fffffffc000,
64'hff7fffff00000081,64'h0001fffffffe0000,64'hfbffffff00000401,64'h000ffffffff00000,
64'hdfffffff00002001,64'h007fffffff800000,64'hfffffffe00010002,64'h03fffffffc000000,
64'hfffffff700080009,64'h1fffffffe0000000,64'hffffffbf00400041,64'hffffffff00000000,
64'hfffffdff02000201,64'hfffffffefffffff9,64'hffffefff10001001,64'hfffffffeffffffc1,
64'hffff7fff80008001,64'hfffffffefffffe01,64'hfffc000300040001,64'hfffffffefffff001,
64'hffe0001f00200001,64'hfffffffeffff8001,64'hff0000ff01000001,64'hfffffffefffc0001,
64'hf80007ff08000001,64'hfffffffeffe00001,64'hc0003fff40000001,64'hfffffffeff000001,
64'h0002000000000002,64'hfffffffef8000001,64'h0010000000000010,64'hfffffffec0000001,
64'h0080000000000080,64'hfffffffd00000001,64'h0400000000000400,64'hffffffef00000001,
64'h2000000000002000,64'hffffff7f00000001,64'h000000010000ffff,64'hfffffbff00000001,
64'h000000080007fff8,64'hffffdfff00000001,64'h00000040003fffc0,64'hfffeffff00000001,
64'h0000020001fffe00,64'hfff7ffff00000001,64'h000010000ffff000,64'hffbfffff00000001,
64'h000080007fff8000,64'hfdffffff00000001,64'h00040003fffc0000,64'hefffffff00000001,
64'h0020001fffe00000,64'h7fffffff00000001,64'h010000ffff000000,64'hfffffffb00000005,
64'h080007fff8000000,64'hffffffdf00000021,64'h40003fffc0000000,64'hfffffeff00000101,
64'h0001fffffffffffe,64'hfffff7ff00000801,64'h000ffffffffffff0,64'hffffbfff00004001,
64'h007fffffffffff80,64'hfffdffff00020001,64'h03fffffffffffc00,64'hffefffff00100001,
64'h1fffffffffffe000,64'hff7fffff00800001,64'h00000000fffeffff,64'hfbffffff04000001
};
  //------------------------
  // 32
  //------------------------
  localparam [2*32-1:0][63:0] NTT_GF64_BWD_WDIV_N32_PHI_L = {
64'hbfffffff40000001,64'h0000000000000002,64'h0000000000000010,64'h0000000000000080,
64'h0000000000000400,64'h0000000000002000,64'h0000000000010000,64'h0000000000080000,
64'h0000000000400000,64'h0000000002000000,64'h0000000010000000,64'h0000000080000000,
64'h0000000400000000,64'h0000002000000000,64'h0000010000000000,64'h0000080000000000,
64'h0000400000000000,64'h0002000000000000,64'h0010000000000000,64'h0080000000000000,
64'h0400000000000000,64'h2000000000000000,64'h00000000ffffffff,64'h00000007fffffff8,
64'h0000003fffffffc0,64'h000001fffffffe00,64'h00000ffffffff000,64'h00007fffffff8000,
64'h0003fffffffc0000,64'h001fffffffe00000,64'h00ffffffff000000,64'h07fffffff8000000,
64'h3fffffffc0000000,64'hfffffffeffffffff,64'hfffffffefffffff1,64'hfffffffeffffff81,
64'hfffffffefffffc01,64'hfffffffeffffe001,64'hfffffffeffff0001,64'hfffffffefff80001,
64'hfffffffeffc00001,64'hfffffffefe000001,64'hfffffffef0000001,64'hfffffffe80000001,
64'hfffffffb00000001,64'hffffffdf00000001,64'hfffffeff00000001,64'hfffff7ff00000001,
64'hffffbfff00000001,64'hfffdffff00000001,64'hffefffff00000001,64'hff7fffff00000001,
64'hfbffffff00000001,64'hdfffffff00000001,64'hfffffffe00000002,64'hfffffff700000009,
64'hffffffbf00000041,64'hfffffdff00000201,64'hffffefff00001001,64'hffff7fff00008001,
64'hfffbffff00040001,64'hffdfffff00200001,64'hfeffffff01000001,64'hf7ffffff08000001
};
  //------------------------
  // 16
  //------------------------
  localparam [2*16-1:0][63:0] NTT_GF64_BWD_WDIV_N16_PHI_L = {
64'h0000000000000004,64'h0000000000000100,64'h0000000000004000,64'h0000000000100000,
64'h0000000004000000,64'h0000000100000000,64'h0000004000000000,64'h0000100000000000,
64'h0004000000000000,64'h0100000000000000,64'h4000000000000000,64'h0000000ffffffff0,
64'h000003fffffffc00,64'h0000ffffffff0000,64'h003fffffffc00000,64'h0ffffffff0000000,
64'hfffffffefffffffd,64'hfffffffeffffff01,64'hfffffffeffffc001,64'hfffffffefff00001,
64'hfffffffefc000001,64'hfffffffe00000001,64'hffffffbf00000001,64'hffffefff00000001,
64'hfffbffff00000001,64'hfeffffff00000001,64'hbfffffff00000001,64'hffffffef00000011,
64'hfffffbff00000401,64'hfffeffff00010001,64'hffbfffff00400001,64'hefffffff10000001
};
  //------------------------
  // 8
  //------------------------
  localparam [2*8-1:0][63:0] NTT_GF64_BWD_WDIV_N8_PHI_L = {
64'h0000000000000200,64'h0000000000200000,64'h0000000200000000,64'h0000200000000000,
64'h0200000000000000,64'h0000001fffffffe0,64'h0001fffffffe0000,64'h1fffffffe0000000,
64'hfffffffefffffe01,64'hfffffffeffe00001,64'hfffffffd00000001,64'hffffdfff00000001,
64'hfdffffff00000001,64'hffffffdf00000021,64'hfffdffff00020001,64'hdfffffff20000001
};
  //------------------------
  // 4
  //------------------------
  localparam [2*4-1:0][63:0] NTT_GF64_BWD_WDIV_N4_PHI_L = {
64'h0000000000400000,64'h0000400000000000,64'h0000003fffffffc0,64'h3fffffffc0000000,
64'hfffffffeffc00001,64'hffffbfff00000001,64'hffffffbf00000041,64'hbfffffff40000001
};

endpackage