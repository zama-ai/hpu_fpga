// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// NTT core (ntt_core) definition package.
// This package defines the key localparams of ntt_core.
// It's content is exported by ntt_core_common_param_pkg.
// Do not use this package directly. Use ntt_core_common_param_pkg.
// ==============================================================================================

package ntt_core_common_div_definition_pkg;
  localparam  int           BWD_PSI_DIV   = 1; // PSI/BWD_PSI_DIV: number of butterflies for INTT
endpackage

