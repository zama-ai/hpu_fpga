// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in any top.
// Should not be used as is.
// Should be imported by top_common_param_pkg.
// ==============================================================================================

package top_common_pc_definition_pkg;
  localparam int PEM_PC  = 1;
  localparam int GLWE_PC = 1;
  localparam int BSK_PC  = 4;
  localparam int KSK_PC  = 4;
endpackage
