// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// bsk_network definition package
// Contains localparams needed for the bsk network.
// ==============================================================================================

package bsk_ntw_common_definition_pkg;
  localparam  int BSK_DIST_COEF_NB          = 48;//64; // should divide BSK_ITER_COEF_NB

endpackage
