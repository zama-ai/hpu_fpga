// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// This file is only a place to set Verilog `define and is only used in simulation
// ==============================================================================================

`ifndef TOP_DEFINES
`define TOP_DEFINES

`define MEMORY_FILE_PATH ""

`endif
