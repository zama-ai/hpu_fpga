// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Parameters that defines the NTT.
// ==============================================================================================

package param_ntt_pkg;
  import param_ntt_definition_pkg::*;

  export param_ntt_definition_pkg::MOD_NTT_W;
  export param_ntt_definition_pkg::MOD_NTT;
  export param_ntt_definition_pkg::MOD_NTT_TYPE;
  export param_ntt_definition_pkg::MOD_NTT_INV_TYPE;
  export param_ntt_definition_pkg::MOD_NTT_NAME;
  export param_ntt_definition_pkg::MOD_NTT_NAME_S;

  // Add here any functions or localparam that are deduced from the previous ones.
endpackage
