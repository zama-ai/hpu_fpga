// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in bsk_manager.
// This package is used to ease the use of several values for these parameters.
// Do not use this package directly. Use bsk_mgr_common_param_pkg.
// ==============================================================================================

package bsk_mgr_common_cut_definition_pkg;
  localparam int BSK_CUT_NB  = 16;
endpackage
