// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in the top.
// Should not be used as is.
// Should be imported by top_common_param_pkg.
// ==============================================================================================

package top_common_top_definition_pkg;
  import common_definition_pkg::*;

  //== Top
  localparam top_name_e        TOP        = TOP_NAME_HPU;

endpackage
