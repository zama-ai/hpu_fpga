// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Package used by ntt_core_gf64_phi.
//
// ==============================================================================================

package ntt_core_gf64_phi_pkg;

// ============================================================================================== //
// Functions
// ============================================================================================== //
  // Reverse <v> in range <range>, in base 2
  // range should be a power of 2
  function [31:0] reverse_int (input [31:0] v, input [31:0] range);
    var [31:0] sz;
    var [31:0] res;

    sz = $clog2(range);
    res = '0;
    for (int i=0; i<32; i=i+1)
      if (i < sz)
        res = res * 2 + v[i];
    return res;
  endfunction


endpackage
