// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in any top.
// Should not be used as is.
// Should be imported by top_common_param_pkg.
// ==============================================================================================

package top_common_pcmax_definition_pkg;
  localparam int PEM_PC_MAX  = 2;
  localparam int GLWE_PC_MAX = 1;
  localparam int BSK_PC_MAX  = 8;
  localparam int KSK_PC_MAX  = 8;
endpackage
