// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// NTT core (ntt_core) definition package.
// This package defines the key localparams of ntt_core.
// It's content is exported by ntt_core_common_param_pkg.
// Do not use this package directly. Use ntt_core_common_param_pkg.
// ==============================================================================================

package ntt_core_common_psi_definition_pkg;
  localparam  int           PSI           = 32; // Number of butterflies
endpackage

