// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  : Common localparams for ucore
// ----------------------------------------------------------------------------------------------
//
// Contain ucore register layout and interface width.
// ==============================================================================================

package ucore_pkg;

  localparam int UCORE_FIFO_DEPTH = 64;
  localparam int ACKQ_RD_ERR = 'hdeadc0de;
endpackage

