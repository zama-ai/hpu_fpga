// ==============================================================================================
// BSD 3-Clause Clear License
// Copyright © 2025 ZAMA. All rights reserved.
// ----------------------------------------------------------------------------------------------
// Description  :
// ----------------------------------------------------------------------------------------------
//
// Definition of localparams used in pep_key_switch.
// ==============================================================================================

package pep_ks_common_definition_pkg;
  // Number of coefficients to be processed in parallel
  localparam int LBY = 16;
  localparam int LBX = 4;
  localparam int LBZ = 3;
endpackage
